magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771281926
<< metal1 >>
rect 576 38576 79584 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 79584 38576
rect 576 38512 79584 38536
rect 64107 38324 64149 38333
rect 64107 38284 64108 38324
rect 64148 38284 64149 38324
rect 64107 38275 64149 38284
rect 58059 38240 58101 38249
rect 58059 38200 58060 38240
rect 58100 38200 58101 38240
rect 58059 38191 58101 38200
rect 58251 38240 58293 38249
rect 58251 38200 58252 38240
rect 58292 38200 58293 38240
rect 58251 38191 58293 38200
rect 58339 38240 58397 38241
rect 58339 38200 58348 38240
rect 58388 38200 58397 38240
rect 58339 38199 58397 38200
rect 59403 38240 59445 38249
rect 59403 38200 59404 38240
rect 59444 38200 59445 38240
rect 59403 38191 59445 38200
rect 63531 38240 63573 38249
rect 63531 38200 63532 38240
rect 63572 38200 63573 38240
rect 63531 38191 63573 38200
rect 63723 38240 63765 38249
rect 63723 38200 63724 38240
rect 63764 38200 63765 38240
rect 63723 38191 63765 38200
rect 63811 38240 63869 38241
rect 63811 38200 63820 38240
rect 63860 38200 63869 38240
rect 63811 38199 63869 38200
rect 64003 38240 64061 38241
rect 64003 38200 64012 38240
rect 64052 38200 64061 38240
rect 64003 38199 64061 38200
rect 64203 38240 64245 38249
rect 64203 38200 64204 38240
rect 64244 38200 64245 38240
rect 64203 38191 64245 38200
rect 67459 38240 67517 38241
rect 67459 38200 67468 38240
rect 67508 38200 67517 38240
rect 67459 38199 67517 38200
rect 68043 38240 68085 38249
rect 68043 38200 68044 38240
rect 68084 38200 68085 38240
rect 68043 38191 68085 38200
rect 68139 38240 68181 38249
rect 68139 38200 68140 38240
rect 68180 38200 68181 38240
rect 68139 38191 68181 38200
rect 68235 38240 68277 38249
rect 68235 38200 68236 38240
rect 68276 38200 68277 38240
rect 68235 38191 68277 38200
rect 68331 38240 68373 38249
rect 68331 38200 68332 38240
rect 68372 38200 68373 38240
rect 68331 38191 68373 38200
rect 68707 38240 68765 38241
rect 68707 38200 68716 38240
rect 68756 38200 68765 38240
rect 68707 38199 68765 38200
rect 68811 38240 68853 38249
rect 68811 38200 68812 38240
rect 68852 38200 68853 38240
rect 68811 38191 68853 38200
rect 69003 38240 69045 38249
rect 69003 38200 69004 38240
rect 69044 38200 69045 38240
rect 69003 38191 69045 38200
rect 70155 38240 70197 38249
rect 70155 38200 70156 38240
rect 70196 38200 70197 38240
rect 70155 38191 70197 38200
rect 71403 38240 71445 38249
rect 71403 38200 71404 38240
rect 71444 38200 71445 38240
rect 71403 38191 71445 38200
rect 72739 38240 72797 38241
rect 72739 38200 72748 38240
rect 72788 38200 72797 38240
rect 72739 38199 72797 38200
rect 76867 38240 76925 38241
rect 76867 38200 76876 38240
rect 76916 38200 76925 38240
rect 76867 38199 76925 38200
rect 77163 38240 77205 38249
rect 77163 38200 77164 38240
rect 77204 38200 77205 38240
rect 77163 38191 77205 38200
rect 77259 38240 77301 38249
rect 77259 38200 77260 38240
rect 77300 38200 77301 38240
rect 77259 38191 77301 38200
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 57283 38156 57341 38157
rect 57283 38116 57292 38156
rect 57332 38116 57341 38156
rect 57283 38115 57341 38116
rect 57667 38156 57725 38157
rect 57667 38116 57676 38156
rect 57716 38116 57725 38156
rect 57667 38115 57725 38116
rect 59971 38156 60029 38157
rect 59971 38116 59980 38156
rect 60020 38116 60029 38156
rect 59971 38115 60029 38116
rect 67843 38156 67901 38157
rect 67843 38116 67852 38156
rect 67892 38116 67901 38156
rect 67843 38115 67901 38116
rect 69387 38156 69429 38165
rect 69387 38116 69388 38156
rect 69428 38116 69429 38156
rect 69387 38107 69429 38116
rect 70635 38156 70677 38165
rect 70635 38116 70636 38156
rect 70676 38116 70677 38156
rect 70635 38107 70677 38116
rect 56427 38072 56469 38081
rect 56427 38032 56428 38072
rect 56468 38032 56469 38072
rect 56427 38023 56469 38032
rect 57867 38072 57909 38081
rect 57867 38032 57868 38072
rect 57908 38032 57909 38072
rect 57867 38023 57909 38032
rect 60171 38072 60213 38081
rect 60171 38032 60172 38072
rect 60212 38032 60213 38072
rect 60171 38023 60213 38032
rect 61899 38072 61941 38081
rect 61899 38032 61900 38072
rect 61940 38032 61941 38072
rect 61899 38023 61941 38032
rect 64587 38072 64629 38081
rect 64587 38032 64588 38072
rect 64628 38032 64629 38072
rect 64587 38023 64629 38032
rect 66219 38072 66261 38081
rect 66219 38032 66220 38072
rect 66260 38032 66261 38072
rect 66219 38023 66261 38032
rect 71979 38072 72021 38081
rect 71979 38032 71980 38072
rect 72020 38032 72021 38072
rect 71979 38023 72021 38032
rect 73995 38072 74037 38081
rect 73995 38032 73996 38072
rect 74036 38032 74037 38072
rect 73995 38023 74037 38032
rect 76011 38072 76053 38081
rect 76011 38032 76012 38072
rect 76052 38032 76053 38072
rect 76011 38023 76053 38032
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 57483 37988 57525 37997
rect 57483 37948 57484 37988
rect 57524 37948 57525 37988
rect 57483 37939 57525 37948
rect 58059 37988 58101 37997
rect 58059 37948 58060 37988
rect 58100 37948 58101 37988
rect 58059 37939 58101 37948
rect 58827 37988 58869 37997
rect 58827 37948 58828 37988
rect 58868 37948 58869 37988
rect 58827 37939 58869 37948
rect 59787 37988 59829 37997
rect 59787 37948 59788 37988
rect 59828 37948 59829 37988
rect 59787 37939 59829 37948
rect 63531 37988 63573 37997
rect 63531 37948 63532 37988
rect 63572 37948 63573 37988
rect 63531 37939 63573 37948
rect 67659 37988 67701 37997
rect 67659 37948 67660 37988
rect 67700 37948 67701 37988
rect 67659 37939 67701 37948
rect 69003 37988 69045 37997
rect 69003 37948 69004 37988
rect 69044 37948 69045 37988
rect 69003 37939 69045 37948
rect 73035 37988 73077 37997
rect 73035 37948 73036 37988
rect 73076 37948 73077 37988
rect 73035 37939 73077 37948
rect 77539 37988 77597 37989
rect 77539 37948 77548 37988
rect 77588 37948 77597 37988
rect 77539 37947 77597 37948
rect 576 37820 79584 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 79584 37820
rect 576 37756 79584 37780
rect 67755 37652 67797 37661
rect 67755 37612 67756 37652
rect 67796 37612 67797 37652
rect 67755 37603 67797 37612
rect 54891 37568 54933 37577
rect 54891 37528 54892 37568
rect 54932 37528 54933 37568
rect 54891 37519 54933 37528
rect 78507 37568 78549 37577
rect 78507 37528 78508 37568
rect 78548 37528 78549 37568
rect 78507 37519 78549 37528
rect 67555 37484 67613 37485
rect 67555 37444 67564 37484
rect 67604 37444 67613 37484
rect 67555 37443 67613 37444
rect 55467 37400 55509 37409
rect 55467 37360 55468 37400
rect 55508 37360 55509 37400
rect 55467 37351 55509 37360
rect 55659 37400 55701 37409
rect 55659 37360 55660 37400
rect 55700 37360 55701 37400
rect 55659 37351 55701 37360
rect 55747 37400 55805 37401
rect 55747 37360 55756 37400
rect 55796 37360 55805 37400
rect 55747 37359 55805 37360
rect 55947 37400 55989 37409
rect 55947 37360 55948 37400
rect 55988 37360 55989 37400
rect 55947 37351 55989 37360
rect 56323 37400 56381 37401
rect 56323 37360 56332 37400
rect 56372 37360 56381 37400
rect 56323 37359 56381 37360
rect 57187 37400 57245 37401
rect 57187 37360 57196 37400
rect 57236 37360 57245 37400
rect 57187 37359 57245 37360
rect 58539 37400 58581 37409
rect 58539 37360 58540 37400
rect 58580 37360 58581 37400
rect 58539 37351 58581 37360
rect 58635 37400 58677 37409
rect 58635 37360 58636 37400
rect 58676 37360 58677 37400
rect 58635 37351 58677 37360
rect 58731 37400 58773 37409
rect 58731 37360 58732 37400
rect 58772 37360 58773 37400
rect 58731 37351 58773 37360
rect 59491 37400 59549 37401
rect 59491 37360 59500 37400
rect 59540 37360 59549 37400
rect 59491 37359 59549 37360
rect 60355 37400 60413 37401
rect 60355 37360 60364 37400
rect 60404 37360 60413 37400
rect 60355 37359 60413 37360
rect 62083 37400 62141 37401
rect 62083 37360 62092 37400
rect 62132 37360 62141 37400
rect 62083 37359 62141 37360
rect 62947 37400 63005 37401
rect 62947 37360 62956 37400
rect 62996 37360 63005 37400
rect 62947 37359 63005 37360
rect 64299 37400 64341 37409
rect 64299 37360 64300 37400
rect 64340 37360 64341 37400
rect 64299 37351 64341 37360
rect 64675 37400 64733 37401
rect 64675 37360 64684 37400
rect 64724 37360 64733 37400
rect 64675 37359 64733 37360
rect 65539 37400 65597 37401
rect 65539 37360 65548 37400
rect 65588 37360 65597 37400
rect 65539 37359 65597 37360
rect 67083 37400 67125 37409
rect 67083 37360 67084 37400
rect 67124 37360 67125 37400
rect 67083 37351 67125 37360
rect 67275 37400 67317 37409
rect 67275 37360 67276 37400
rect 67316 37360 67317 37400
rect 67275 37351 67317 37360
rect 67363 37400 67421 37401
rect 67363 37360 67372 37400
rect 67412 37360 67421 37400
rect 67363 37359 67421 37360
rect 68035 37400 68093 37401
rect 68035 37360 68044 37400
rect 68084 37360 68093 37400
rect 68035 37359 68093 37360
rect 68331 37400 68373 37409
rect 68331 37360 68332 37400
rect 68372 37360 68373 37400
rect 68331 37351 68373 37360
rect 69099 37400 69141 37409
rect 69099 37360 69100 37400
rect 69140 37360 69141 37400
rect 69099 37351 69141 37360
rect 69475 37400 69533 37401
rect 69475 37360 69484 37400
rect 69524 37360 69533 37400
rect 69475 37359 69533 37360
rect 70339 37400 70397 37401
rect 70339 37360 70348 37400
rect 70388 37360 70397 37400
rect 70339 37359 70397 37360
rect 72747 37400 72789 37409
rect 72747 37360 72748 37400
rect 72788 37360 72789 37400
rect 72747 37351 72789 37360
rect 72843 37400 72885 37409
rect 72843 37360 72844 37400
rect 72884 37360 72885 37400
rect 72843 37351 72885 37360
rect 72939 37400 72981 37409
rect 72939 37360 72940 37400
rect 72980 37360 72981 37400
rect 72939 37351 72981 37360
rect 73227 37400 73269 37409
rect 73227 37360 73228 37400
rect 73268 37360 73269 37400
rect 73507 37400 73565 37401
rect 73227 37351 73269 37360
rect 73419 37358 73461 37367
rect 73507 37360 73516 37400
rect 73556 37360 73565 37400
rect 73507 37359 73565 37360
rect 73707 37400 73749 37409
rect 73707 37360 73708 37400
rect 73748 37360 73749 37400
rect 59115 37316 59157 37325
rect 59115 37276 59116 37316
rect 59156 37276 59157 37316
rect 59115 37267 59157 37276
rect 61707 37316 61749 37325
rect 61707 37276 61708 37316
rect 61748 37276 61749 37316
rect 61707 37267 61749 37276
rect 68427 37316 68469 37325
rect 68427 37276 68428 37316
rect 68468 37276 68469 37316
rect 68427 37267 68469 37276
rect 73035 37316 73077 37325
rect 73035 37276 73036 37316
rect 73076 37276 73077 37316
rect 73419 37318 73420 37358
rect 73460 37318 73461 37358
rect 73707 37351 73749 37360
rect 73899 37400 73941 37409
rect 73899 37360 73900 37400
rect 73940 37360 73941 37400
rect 73899 37351 73941 37360
rect 73987 37400 74045 37401
rect 73987 37360 73996 37400
rect 74036 37360 74045 37400
rect 73987 37359 74045 37360
rect 74283 37400 74325 37409
rect 74283 37360 74284 37400
rect 74324 37360 74325 37400
rect 74283 37351 74325 37360
rect 74475 37400 74517 37409
rect 74475 37360 74476 37400
rect 74516 37360 74517 37400
rect 74475 37351 74517 37360
rect 74563 37400 74621 37401
rect 74563 37360 74572 37400
rect 74612 37360 74621 37400
rect 74563 37359 74621 37360
rect 75051 37400 75093 37409
rect 75051 37360 75052 37400
rect 75092 37360 75093 37400
rect 75051 37351 75093 37360
rect 75147 37400 75189 37409
rect 75147 37360 75148 37400
rect 75188 37360 75189 37400
rect 75147 37351 75189 37360
rect 75243 37400 75285 37409
rect 75243 37360 75244 37400
rect 75284 37360 75285 37400
rect 75243 37351 75285 37360
rect 75907 37400 75965 37401
rect 75907 37360 75916 37400
rect 75956 37360 75965 37400
rect 75907 37359 75965 37360
rect 76771 37400 76829 37401
rect 76771 37360 76780 37400
rect 76820 37360 76829 37400
rect 76771 37359 76829 37360
rect 78115 37400 78173 37401
rect 78115 37360 78124 37400
rect 78164 37360 78173 37400
rect 78115 37359 78173 37360
rect 78315 37400 78357 37409
rect 78315 37360 78316 37400
rect 78356 37360 78357 37400
rect 78315 37351 78357 37360
rect 73419 37309 73461 37318
rect 74379 37316 74421 37325
rect 73035 37267 73077 37276
rect 74379 37276 74380 37316
rect 74420 37276 74421 37316
rect 74379 37267 74421 37276
rect 75531 37316 75573 37325
rect 75531 37276 75532 37316
rect 75572 37276 75573 37316
rect 75531 37267 75573 37276
rect 78219 37316 78261 37325
rect 78219 37276 78220 37316
rect 78260 37276 78261 37316
rect 78219 37267 78261 37276
rect 55555 37232 55613 37233
rect 55555 37192 55564 37232
rect 55604 37192 55613 37232
rect 55555 37191 55613 37192
rect 58339 37232 58397 37233
rect 58339 37192 58348 37232
rect 58388 37192 58397 37232
rect 58339 37191 58397 37192
rect 58819 37232 58877 37233
rect 58819 37192 58828 37232
rect 58868 37192 58877 37232
rect 58819 37191 58877 37192
rect 61507 37232 61565 37233
rect 61507 37192 61516 37232
rect 61556 37192 61565 37232
rect 61507 37191 61565 37192
rect 64099 37232 64157 37233
rect 64099 37192 64108 37232
rect 64148 37192 64157 37232
rect 64099 37191 64157 37192
rect 66691 37232 66749 37233
rect 66691 37192 66700 37232
rect 66740 37192 66749 37232
rect 66691 37191 66749 37192
rect 67171 37232 67229 37233
rect 67171 37192 67180 37232
rect 67220 37192 67229 37232
rect 67171 37191 67229 37192
rect 67755 37232 67797 37241
rect 67755 37192 67756 37232
rect 67796 37192 67797 37232
rect 71491 37232 71549 37233
rect 67755 37183 67797 37192
rect 68715 37190 68757 37199
rect 71491 37192 71500 37232
rect 71540 37192 71549 37232
rect 71491 37191 71549 37192
rect 73315 37232 73373 37233
rect 73315 37192 73324 37232
rect 73364 37192 73373 37232
rect 73315 37191 73373 37192
rect 73795 37232 73853 37233
rect 73795 37192 73804 37232
rect 73844 37192 73853 37232
rect 73795 37191 73853 37192
rect 75331 37232 75389 37233
rect 75331 37192 75340 37232
rect 75380 37192 75389 37232
rect 75331 37191 75389 37192
rect 77923 37232 77981 37233
rect 77923 37192 77932 37232
rect 77972 37192 77981 37232
rect 77923 37191 77981 37192
rect 68715 37150 68716 37190
rect 68756 37150 68757 37190
rect 68715 37141 68757 37150
rect 576 37064 79584 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 79584 37064
rect 576 37000 79584 37024
rect 57091 36896 57149 36897
rect 57091 36856 57100 36896
rect 57140 36856 57149 36896
rect 57091 36855 57149 36856
rect 59203 36896 59261 36897
rect 59203 36856 59212 36896
rect 59252 36856 59261 36896
rect 59203 36855 59261 36856
rect 60259 36896 60317 36897
rect 60259 36856 60268 36896
rect 60308 36856 60317 36896
rect 60259 36855 60317 36856
rect 61987 36896 62045 36897
rect 61987 36856 61996 36896
rect 62036 36856 62045 36896
rect 61987 36855 62045 36856
rect 68131 36896 68189 36897
rect 68131 36856 68140 36896
rect 68180 36856 68189 36896
rect 68131 36855 68189 36856
rect 76195 36896 76253 36897
rect 76195 36856 76204 36896
rect 76244 36856 76253 36896
rect 76195 36855 76253 36856
rect 79459 36896 79517 36897
rect 79459 36856 79468 36896
rect 79508 36856 79517 36896
rect 79459 36855 79517 36856
rect 54411 36812 54453 36821
rect 54411 36772 54412 36812
rect 54452 36772 54453 36812
rect 54411 36763 54453 36772
rect 59691 36812 59733 36821
rect 59691 36772 59692 36812
rect 59732 36772 59733 36812
rect 59691 36763 59733 36772
rect 63531 36812 63573 36821
rect 63531 36772 63532 36812
rect 63572 36772 63573 36812
rect 63531 36763 63573 36772
rect 69003 36812 69045 36821
rect 69003 36772 69004 36812
rect 69044 36772 69045 36812
rect 69003 36763 69045 36772
rect 69387 36812 69429 36821
rect 69387 36772 69388 36812
rect 69428 36772 69429 36812
rect 69387 36763 69429 36772
rect 73323 36812 73365 36821
rect 73323 36772 73324 36812
rect 73364 36772 73365 36812
rect 73323 36763 73365 36772
rect 73515 36812 73557 36821
rect 73515 36772 73516 36812
rect 73556 36772 73557 36812
rect 73515 36763 73557 36772
rect 54787 36728 54845 36729
rect 54787 36688 54796 36728
rect 54836 36688 54845 36728
rect 54787 36687 54845 36688
rect 55651 36728 55709 36729
rect 55651 36688 55660 36728
rect 55700 36688 55709 36728
rect 55651 36687 55709 36688
rect 57003 36728 57045 36737
rect 57003 36688 57004 36728
rect 57044 36688 57045 36728
rect 57003 36679 57045 36688
rect 57195 36728 57237 36737
rect 57195 36688 57196 36728
rect 57236 36688 57237 36728
rect 57195 36679 57237 36688
rect 57283 36728 57341 36729
rect 57283 36688 57292 36728
rect 57332 36688 57341 36728
rect 57283 36687 57341 36688
rect 58243 36728 58301 36729
rect 58243 36688 58252 36728
rect 58292 36688 58301 36728
rect 58243 36687 58301 36688
rect 58539 36728 58581 36737
rect 58539 36688 58540 36728
rect 58580 36688 58581 36728
rect 58539 36679 58581 36688
rect 58635 36728 58677 36737
rect 58635 36688 58636 36728
rect 58676 36688 58677 36728
rect 58635 36679 58677 36688
rect 59115 36728 59157 36737
rect 59115 36688 59116 36728
rect 59156 36688 59157 36728
rect 59115 36679 59157 36688
rect 59307 36728 59349 36737
rect 59307 36688 59308 36728
rect 59348 36688 59349 36728
rect 59307 36679 59349 36688
rect 59395 36728 59453 36729
rect 59395 36688 59404 36728
rect 59444 36688 59453 36728
rect 59395 36687 59453 36688
rect 59587 36728 59645 36729
rect 59587 36688 59596 36728
rect 59636 36688 59645 36728
rect 59587 36687 59645 36688
rect 59787 36728 59829 36737
rect 59787 36688 59788 36728
rect 59828 36688 59829 36728
rect 59787 36679 59829 36688
rect 60171 36728 60213 36737
rect 60171 36688 60172 36728
rect 60212 36688 60213 36728
rect 60171 36679 60213 36688
rect 60363 36728 60405 36737
rect 60363 36688 60364 36728
rect 60404 36688 60405 36728
rect 60363 36679 60405 36688
rect 60451 36728 60509 36729
rect 60451 36688 60460 36728
rect 60500 36688 60509 36728
rect 60451 36687 60509 36688
rect 61419 36728 61461 36737
rect 61419 36688 61420 36728
rect 61460 36688 61461 36728
rect 61419 36679 61461 36688
rect 61515 36728 61557 36737
rect 61515 36688 61516 36728
rect 61556 36688 61557 36728
rect 61515 36679 61557 36688
rect 61611 36728 61653 36737
rect 61611 36688 61612 36728
rect 61652 36688 61653 36728
rect 61611 36679 61653 36688
rect 61707 36728 61749 36737
rect 61707 36688 61708 36728
rect 61748 36688 61749 36728
rect 61707 36679 61749 36688
rect 61899 36728 61941 36737
rect 61899 36688 61900 36728
rect 61940 36688 61941 36728
rect 61899 36679 61941 36688
rect 62091 36728 62133 36737
rect 62091 36688 62092 36728
rect 62132 36688 62133 36728
rect 62091 36679 62133 36688
rect 62179 36728 62237 36729
rect 62179 36688 62188 36728
rect 62228 36688 62237 36728
rect 62179 36687 62237 36688
rect 63139 36728 63197 36729
rect 63139 36688 63148 36728
rect 63188 36688 63197 36728
rect 63139 36687 63197 36688
rect 63435 36728 63477 36737
rect 63435 36688 63436 36728
rect 63476 36688 63477 36728
rect 63435 36679 63477 36688
rect 64011 36728 64053 36737
rect 64011 36688 64012 36728
rect 64052 36688 64053 36728
rect 64011 36679 64053 36688
rect 64195 36728 64253 36729
rect 64195 36688 64204 36728
rect 64244 36688 64253 36728
rect 64195 36687 64253 36688
rect 65739 36728 65781 36737
rect 65739 36688 65740 36728
rect 65780 36688 65781 36728
rect 65739 36679 65781 36688
rect 66115 36728 66173 36729
rect 66115 36688 66124 36728
rect 66164 36688 66173 36728
rect 66115 36687 66173 36688
rect 66979 36728 67037 36729
rect 66979 36688 66988 36728
rect 67028 36688 67037 36728
rect 66979 36687 67037 36688
rect 68427 36728 68469 36737
rect 68427 36688 68428 36728
rect 68468 36688 68469 36728
rect 68427 36679 68469 36688
rect 68619 36728 68661 36737
rect 68619 36688 68620 36728
rect 68660 36688 68661 36728
rect 68619 36679 68661 36688
rect 68707 36728 68765 36729
rect 68707 36688 68716 36728
rect 68756 36688 68765 36728
rect 68707 36687 68765 36688
rect 68907 36728 68949 36737
rect 68907 36688 68908 36728
rect 68948 36688 68949 36728
rect 69283 36728 69341 36729
rect 68907 36679 68949 36688
rect 69086 36705 69144 36706
rect 69086 36665 69095 36705
rect 69135 36665 69144 36705
rect 69283 36688 69292 36728
rect 69332 36688 69341 36728
rect 69283 36687 69341 36688
rect 69483 36728 69525 36737
rect 69483 36688 69484 36728
rect 69524 36688 69525 36728
rect 69483 36679 69525 36688
rect 72067 36728 72125 36729
rect 72067 36688 72076 36728
rect 72116 36688 72125 36728
rect 72067 36687 72125 36688
rect 72931 36728 72989 36729
rect 72931 36688 72940 36728
rect 72980 36688 72989 36728
rect 72931 36687 72989 36688
rect 73891 36728 73949 36729
rect 73891 36688 73900 36728
rect 73940 36688 73949 36728
rect 73891 36687 73949 36688
rect 74755 36728 74813 36729
rect 74755 36688 74764 36728
rect 74804 36688 74813 36728
rect 74755 36687 74813 36688
rect 76107 36728 76149 36737
rect 76107 36688 76108 36728
rect 76148 36688 76149 36728
rect 76107 36679 76149 36688
rect 76299 36728 76341 36737
rect 76299 36688 76300 36728
rect 76340 36688 76341 36728
rect 76299 36679 76341 36688
rect 76387 36728 76445 36729
rect 76387 36688 76396 36728
rect 76436 36688 76445 36728
rect 76387 36687 76445 36688
rect 76587 36728 76629 36737
rect 76587 36688 76588 36728
rect 76628 36688 76629 36728
rect 76587 36679 76629 36688
rect 76779 36728 76821 36737
rect 76779 36688 76780 36728
rect 76820 36688 76821 36728
rect 76779 36679 76821 36688
rect 76867 36728 76925 36729
rect 76867 36688 76876 36728
rect 76916 36688 76925 36728
rect 76867 36687 76925 36688
rect 77067 36728 77109 36737
rect 77067 36688 77068 36728
rect 77108 36688 77109 36728
rect 77067 36679 77109 36688
rect 77443 36728 77501 36729
rect 77443 36688 77452 36728
rect 77492 36688 77501 36728
rect 77443 36687 77501 36688
rect 78307 36728 78365 36729
rect 78307 36688 78316 36728
rect 78356 36688 78365 36728
rect 78307 36687 78365 36688
rect 69086 36664 69144 36665
rect 63811 36560 63869 36561
rect 63811 36520 63820 36560
rect 63860 36520 63869 36560
rect 63811 36519 63869 36520
rect 64107 36560 64149 36569
rect 64107 36520 64108 36560
rect 64148 36520 64149 36560
rect 64107 36511 64149 36520
rect 69675 36560 69717 36569
rect 69675 36520 69676 36560
rect 69716 36520 69717 36560
rect 69675 36511 69717 36520
rect 76587 36560 76629 36569
rect 76587 36520 76588 36560
rect 76628 36520 76629 36560
rect 76587 36511 76629 36520
rect 56803 36476 56861 36477
rect 56803 36436 56812 36476
rect 56852 36436 56861 36476
rect 56803 36435 56861 36436
rect 58915 36476 58973 36477
rect 58915 36436 58924 36476
rect 58964 36436 58973 36476
rect 58915 36435 58973 36436
rect 68427 36476 68469 36485
rect 68427 36436 68428 36476
rect 68468 36436 68469 36476
rect 68427 36427 68469 36436
rect 70915 36476 70973 36477
rect 70915 36436 70924 36476
rect 70964 36436 70973 36476
rect 70915 36435 70973 36436
rect 75907 36476 75965 36477
rect 75907 36436 75916 36476
rect 75956 36436 75965 36476
rect 75907 36435 75965 36436
rect 576 36308 79584 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 79584 36308
rect 576 36244 79584 36268
rect 73707 36140 73749 36149
rect 73707 36100 73708 36140
rect 73748 36100 73749 36140
rect 73707 36091 73749 36100
rect 74091 36140 74133 36149
rect 74091 36100 74092 36140
rect 74132 36100 74133 36140
rect 74091 36091 74133 36100
rect 76491 36140 76533 36149
rect 76491 36100 76492 36140
rect 76532 36100 76533 36140
rect 76491 36091 76533 36100
rect 77547 36140 77589 36149
rect 77547 36100 77548 36140
rect 77588 36100 77589 36140
rect 77547 36091 77589 36100
rect 49131 36056 49173 36065
rect 49131 36016 49132 36056
rect 49172 36016 49173 36056
rect 49131 36007 49173 36016
rect 60267 36056 60309 36065
rect 60267 36016 60268 36056
rect 60308 36016 60309 36056
rect 60267 36007 60309 36016
rect 69483 36056 69525 36065
rect 69483 36016 69484 36056
rect 69524 36016 69525 36056
rect 69483 36007 69525 36016
rect 74667 36056 74709 36065
rect 74667 36016 74668 36056
rect 74708 36016 74709 36056
rect 73411 36014 73469 36015
rect 50947 35972 51005 35973
rect 50947 35932 50956 35972
rect 50996 35932 51005 35972
rect 50947 35931 51005 35932
rect 56803 35972 56861 35973
rect 56803 35932 56812 35972
rect 56852 35932 56861 35972
rect 56803 35931 56861 35932
rect 58923 35972 58965 35981
rect 73411 35974 73420 36014
rect 73460 35974 73469 36014
rect 74667 36007 74709 36016
rect 77835 36056 77877 36065
rect 77835 36016 77836 36056
rect 77876 36016 77877 36056
rect 77835 36007 77877 36016
rect 73411 35973 73469 35974
rect 58923 35932 58924 35972
rect 58964 35932 58965 35972
rect 58923 35923 58965 35932
rect 51243 35888 51285 35897
rect 51243 35848 51244 35888
rect 51284 35848 51285 35888
rect 51243 35839 51285 35848
rect 51427 35888 51485 35889
rect 51427 35848 51436 35888
rect 51476 35848 51485 35888
rect 51427 35847 51485 35848
rect 52387 35888 52445 35889
rect 52387 35848 52396 35888
rect 52436 35848 52445 35888
rect 55755 35888 55797 35897
rect 52387 35847 52445 35848
rect 53251 35877 53309 35878
rect 53251 35837 53260 35877
rect 53300 35837 53309 35877
rect 55755 35848 55756 35888
rect 55796 35848 55797 35888
rect 55755 35839 55797 35848
rect 55851 35888 55893 35897
rect 55851 35848 55852 35888
rect 55892 35848 55893 35888
rect 55851 35839 55893 35848
rect 55947 35888 55989 35897
rect 55947 35848 55948 35888
rect 55988 35848 55989 35888
rect 55947 35839 55989 35848
rect 56043 35888 56085 35897
rect 56043 35848 56044 35888
rect 56084 35848 56085 35888
rect 56043 35839 56085 35848
rect 56227 35888 56285 35889
rect 56227 35848 56236 35888
rect 56276 35848 56285 35888
rect 56227 35847 56285 35848
rect 56427 35888 56469 35897
rect 56427 35848 56428 35888
rect 56468 35848 56469 35888
rect 56427 35839 56469 35848
rect 58827 35888 58869 35897
rect 58827 35848 58828 35888
rect 58868 35848 58869 35888
rect 58827 35839 58869 35848
rect 59011 35888 59069 35889
rect 59011 35848 59020 35888
rect 59060 35848 59069 35888
rect 59011 35847 59069 35848
rect 61323 35888 61365 35897
rect 61323 35848 61324 35888
rect 61364 35848 61365 35888
rect 61323 35839 61365 35848
rect 61515 35888 61557 35897
rect 61515 35848 61516 35888
rect 61556 35848 61557 35888
rect 61515 35839 61557 35848
rect 61603 35888 61661 35889
rect 61603 35848 61612 35888
rect 61652 35848 61661 35888
rect 61603 35847 61661 35848
rect 61899 35888 61941 35897
rect 61899 35848 61900 35888
rect 61940 35848 61941 35888
rect 61899 35839 61941 35848
rect 61995 35888 62037 35897
rect 61995 35848 61996 35888
rect 62036 35848 62037 35888
rect 61995 35839 62037 35848
rect 62091 35888 62133 35897
rect 62091 35848 62092 35888
rect 62132 35848 62133 35888
rect 62091 35839 62133 35848
rect 64579 35888 64637 35889
rect 64579 35848 64588 35888
rect 64628 35848 64637 35888
rect 64579 35847 64637 35848
rect 65443 35888 65501 35889
rect 65443 35848 65452 35888
rect 65492 35848 65501 35888
rect 65443 35847 65501 35848
rect 66795 35888 66837 35897
rect 66795 35848 66796 35888
rect 66836 35848 66837 35888
rect 66795 35839 66837 35848
rect 66987 35888 67029 35897
rect 66987 35848 66988 35888
rect 67028 35848 67029 35888
rect 66987 35839 67029 35848
rect 67075 35888 67133 35889
rect 67075 35848 67084 35888
rect 67124 35848 67133 35888
rect 67075 35847 67133 35848
rect 67267 35888 67325 35889
rect 67267 35848 67276 35888
rect 67316 35848 67325 35888
rect 67267 35847 67325 35848
rect 67371 35888 67413 35897
rect 67371 35848 67372 35888
rect 67412 35848 67413 35888
rect 67371 35839 67413 35848
rect 67467 35888 67509 35897
rect 67467 35848 67468 35888
rect 67508 35848 67509 35888
rect 67467 35839 67509 35848
rect 69675 35888 69717 35897
rect 69675 35848 69676 35888
rect 69716 35848 69717 35888
rect 69675 35839 69717 35848
rect 69867 35888 69909 35897
rect 69867 35848 69868 35888
rect 69908 35848 69909 35888
rect 69867 35839 69909 35848
rect 69955 35888 70013 35889
rect 69955 35848 69964 35888
rect 70004 35848 70013 35888
rect 69955 35847 70013 35848
rect 71883 35888 71925 35897
rect 71883 35848 71884 35888
rect 71924 35848 71925 35888
rect 72163 35888 72221 35889
rect 71883 35839 71925 35848
rect 72075 35874 72117 35883
rect 53251 35836 53309 35837
rect 72075 35834 72076 35874
rect 72116 35834 72117 35874
rect 72163 35848 72172 35888
rect 72212 35848 72221 35888
rect 72163 35847 72221 35848
rect 72739 35888 72797 35889
rect 72739 35848 72748 35888
rect 72788 35848 72797 35888
rect 72739 35847 72797 35848
rect 73035 35888 73077 35897
rect 73035 35848 73036 35888
rect 73076 35848 73077 35888
rect 73035 35839 73077 35848
rect 73603 35888 73661 35889
rect 73603 35848 73612 35888
rect 73652 35848 73661 35888
rect 73603 35847 73661 35848
rect 73803 35888 73845 35897
rect 73803 35848 73804 35888
rect 73844 35848 73845 35888
rect 73803 35839 73845 35848
rect 73995 35888 74037 35897
rect 73995 35848 73996 35888
rect 74036 35848 74037 35888
rect 73995 35839 74037 35848
rect 74179 35888 74237 35889
rect 74179 35848 74188 35888
rect 74228 35848 74237 35888
rect 74179 35847 74237 35848
rect 76107 35888 76149 35897
rect 76107 35848 76108 35888
rect 76148 35848 76149 35888
rect 76107 35839 76149 35848
rect 76203 35888 76245 35897
rect 76203 35848 76204 35888
rect 76244 35848 76245 35888
rect 76203 35839 76245 35848
rect 76299 35888 76341 35897
rect 76299 35848 76300 35888
rect 76340 35848 76341 35888
rect 76299 35839 76341 35848
rect 76491 35888 76533 35897
rect 76491 35848 76492 35888
rect 76532 35848 76533 35888
rect 76491 35839 76533 35848
rect 76683 35888 76725 35897
rect 76683 35848 76684 35888
rect 76724 35848 76725 35888
rect 76683 35839 76725 35848
rect 76771 35888 76829 35889
rect 76771 35848 76780 35888
rect 76820 35848 76829 35888
rect 76771 35847 76829 35848
rect 77059 35888 77117 35889
rect 77059 35848 77068 35888
rect 77108 35848 77117 35888
rect 77059 35847 77117 35848
rect 77259 35888 77301 35897
rect 77259 35848 77260 35888
rect 77300 35848 77301 35888
rect 77259 35839 77301 35848
rect 77443 35888 77501 35889
rect 77443 35848 77452 35888
rect 77492 35848 77501 35888
rect 77443 35847 77501 35848
rect 77643 35888 77685 35897
rect 77643 35848 77644 35888
rect 77684 35848 77685 35888
rect 77643 35839 77685 35848
rect 72075 35825 72117 35834
rect 51339 35804 51381 35813
rect 51339 35764 51340 35804
rect 51380 35764 51381 35804
rect 51339 35755 51381 35764
rect 52011 35804 52053 35813
rect 52011 35764 52012 35804
rect 52052 35764 52053 35804
rect 52011 35755 52053 35764
rect 56331 35804 56373 35813
rect 56331 35764 56332 35804
rect 56372 35764 56373 35804
rect 56331 35755 56373 35764
rect 61419 35804 61461 35813
rect 61419 35764 61420 35804
rect 61460 35764 61461 35804
rect 61419 35755 61461 35764
rect 64203 35804 64245 35813
rect 64203 35764 64204 35804
rect 64244 35764 64245 35804
rect 64203 35755 64245 35764
rect 66891 35804 66933 35813
rect 66891 35764 66892 35804
rect 66932 35764 66933 35804
rect 66891 35755 66933 35764
rect 69771 35804 69813 35813
rect 69771 35764 69772 35804
rect 69812 35764 69813 35804
rect 69771 35755 69813 35764
rect 73131 35804 73173 35813
rect 73131 35764 73132 35804
rect 73172 35764 73173 35804
rect 73131 35755 73173 35764
rect 77163 35804 77205 35813
rect 77163 35764 77164 35804
rect 77204 35764 77205 35804
rect 77163 35755 77205 35764
rect 50763 35720 50805 35729
rect 50763 35680 50764 35720
rect 50804 35680 50805 35720
rect 50763 35671 50805 35680
rect 54403 35720 54461 35721
rect 54403 35680 54412 35720
rect 54452 35680 54461 35720
rect 54403 35679 54461 35680
rect 56619 35720 56661 35729
rect 56619 35680 56620 35720
rect 56660 35680 56661 35720
rect 56619 35671 56661 35680
rect 61795 35720 61853 35721
rect 61795 35680 61804 35720
rect 61844 35680 61853 35720
rect 61795 35679 61853 35680
rect 66595 35720 66653 35721
rect 66595 35680 66604 35720
rect 66644 35680 66653 35720
rect 66595 35679 66653 35680
rect 71971 35720 72029 35721
rect 71971 35680 71980 35720
rect 72020 35680 72029 35720
rect 71971 35679 72029 35680
rect 76003 35720 76061 35721
rect 76003 35680 76012 35720
rect 76052 35680 76061 35720
rect 76003 35679 76061 35680
rect 576 35552 79584 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 79584 35552
rect 576 35488 79584 35512
rect 55171 35384 55229 35385
rect 55171 35344 55180 35384
rect 55220 35344 55229 35384
rect 55171 35343 55229 35344
rect 65827 35384 65885 35385
rect 65827 35344 65836 35384
rect 65876 35344 65885 35384
rect 65827 35343 65885 35344
rect 54795 35300 54837 35309
rect 54795 35260 54796 35300
rect 54836 35260 54837 35300
rect 54795 35251 54837 35260
rect 55563 35300 55605 35309
rect 55563 35260 55564 35300
rect 55604 35260 55605 35300
rect 55563 35251 55605 35260
rect 62667 35300 62709 35309
rect 62667 35260 62668 35300
rect 62708 35260 62709 35300
rect 62667 35251 62709 35260
rect 71403 35300 71445 35309
rect 71403 35260 71404 35300
rect 71444 35260 71445 35300
rect 71403 35251 71445 35260
rect 46539 35216 46581 35225
rect 46539 35176 46540 35216
rect 46580 35176 46581 35216
rect 46539 35167 46581 35176
rect 46731 35216 46773 35225
rect 46731 35176 46732 35216
rect 46772 35176 46773 35216
rect 46731 35167 46773 35176
rect 46819 35216 46877 35217
rect 46819 35176 46828 35216
rect 46868 35176 46877 35216
rect 46819 35175 46877 35176
rect 49603 35216 49661 35217
rect 49603 35176 49612 35216
rect 49652 35176 49661 35216
rect 49603 35175 49661 35176
rect 50467 35216 50525 35217
rect 50467 35176 50476 35216
rect 50516 35176 50525 35216
rect 50467 35175 50525 35176
rect 50859 35216 50901 35225
rect 50859 35176 50860 35216
rect 50900 35176 50901 35216
rect 50859 35167 50901 35176
rect 51339 35216 51381 35225
rect 51339 35176 51340 35216
rect 51380 35176 51381 35216
rect 51339 35167 51381 35176
rect 51435 35216 51477 35225
rect 51435 35176 51436 35216
rect 51476 35176 51477 35216
rect 51435 35167 51477 35176
rect 51715 35216 51773 35217
rect 51715 35176 51724 35216
rect 51764 35176 51773 35216
rect 51715 35175 51773 35176
rect 52003 35216 52061 35217
rect 52003 35176 52012 35216
rect 52052 35176 52061 35216
rect 52299 35216 52341 35225
rect 52003 35175 52061 35176
rect 52099 35202 52157 35203
rect 52099 35162 52108 35202
rect 52148 35162 52157 35202
rect 52299 35176 52300 35216
rect 52340 35176 52341 35216
rect 52299 35167 52341 35176
rect 54691 35216 54749 35217
rect 54691 35176 54700 35216
rect 54740 35176 54749 35216
rect 54691 35175 54749 35176
rect 54891 35216 54933 35225
rect 54891 35176 54892 35216
rect 54932 35176 54933 35216
rect 54891 35167 54933 35176
rect 55083 35216 55125 35225
rect 55083 35176 55084 35216
rect 55124 35176 55125 35216
rect 55083 35167 55125 35176
rect 55275 35216 55317 35225
rect 55275 35176 55276 35216
rect 55316 35176 55317 35216
rect 55939 35216 55997 35217
rect 55275 35167 55317 35176
rect 55389 35205 55431 35214
rect 52099 35161 52157 35162
rect 55389 35165 55390 35205
rect 55430 35165 55431 35205
rect 55939 35176 55948 35216
rect 55988 35176 55997 35216
rect 55939 35175 55997 35176
rect 56803 35216 56861 35217
rect 56803 35176 56812 35216
rect 56852 35176 56861 35216
rect 56803 35175 56861 35176
rect 58155 35216 58197 35225
rect 58155 35176 58156 35216
rect 58196 35176 58197 35216
rect 58155 35167 58197 35176
rect 58347 35216 58389 35225
rect 58347 35176 58348 35216
rect 58388 35176 58389 35216
rect 58347 35167 58389 35176
rect 58435 35216 58493 35217
rect 58435 35176 58444 35216
rect 58484 35176 58493 35216
rect 58435 35175 58493 35176
rect 59787 35216 59829 35225
rect 59787 35176 59788 35216
rect 59828 35176 59829 35216
rect 59787 35167 59829 35176
rect 60163 35216 60221 35217
rect 60163 35176 60172 35216
rect 60212 35176 60221 35216
rect 60163 35175 60221 35176
rect 61027 35216 61085 35217
rect 61027 35176 61036 35216
rect 61076 35176 61085 35216
rect 61027 35175 61085 35176
rect 62763 35216 62805 35225
rect 62763 35176 62764 35216
rect 62804 35176 62805 35216
rect 62763 35167 62805 35176
rect 63043 35216 63101 35217
rect 63043 35176 63052 35216
rect 63092 35176 63101 35216
rect 63043 35175 63101 35176
rect 65931 35216 65973 35225
rect 65931 35176 65932 35216
rect 65972 35176 65973 35216
rect 65931 35167 65973 35176
rect 66027 35216 66069 35225
rect 66027 35176 66028 35216
rect 66068 35176 66069 35216
rect 66027 35167 66069 35176
rect 66123 35216 66165 35225
rect 66123 35176 66124 35216
rect 66164 35176 66165 35216
rect 66123 35167 66165 35176
rect 66403 35216 66461 35217
rect 66403 35176 66412 35216
rect 66452 35176 66461 35216
rect 66403 35175 66461 35176
rect 66699 35216 66741 35225
rect 66699 35176 66700 35216
rect 66740 35176 66741 35216
rect 66699 35167 66741 35176
rect 66795 35216 66837 35225
rect 66795 35176 66796 35216
rect 66836 35176 66837 35216
rect 66795 35167 66837 35176
rect 67467 35216 67509 35225
rect 67467 35176 67468 35216
rect 67508 35176 67509 35216
rect 67467 35167 67509 35176
rect 67843 35216 67901 35217
rect 67843 35176 67852 35216
rect 67892 35176 67901 35216
rect 67843 35175 67901 35176
rect 68707 35216 68765 35217
rect 68707 35176 68716 35216
rect 68756 35176 68765 35216
rect 68707 35175 68765 35176
rect 70443 35216 70485 35225
rect 70443 35176 70444 35216
rect 70484 35176 70485 35216
rect 70443 35167 70485 35176
rect 70539 35216 70581 35225
rect 70539 35176 70540 35216
rect 70580 35176 70581 35216
rect 70539 35167 70581 35176
rect 70635 35216 70677 35225
rect 70635 35176 70636 35216
rect 70676 35176 70677 35216
rect 70635 35167 70677 35176
rect 70731 35216 70773 35225
rect 70731 35176 70732 35216
rect 70772 35176 70773 35216
rect 70731 35167 70773 35176
rect 71011 35216 71069 35217
rect 71011 35176 71020 35216
rect 71060 35176 71069 35216
rect 71011 35175 71069 35176
rect 71307 35216 71349 35225
rect 71307 35176 71308 35216
rect 71348 35176 71349 35216
rect 71307 35167 71349 35176
rect 71883 35216 71925 35225
rect 71883 35176 71884 35216
rect 71924 35176 71925 35216
rect 71883 35167 71925 35176
rect 72075 35216 72117 35225
rect 72075 35176 72076 35216
rect 72116 35176 72117 35216
rect 72075 35167 72117 35176
rect 72163 35216 72221 35217
rect 72163 35176 72172 35216
rect 72212 35176 72221 35216
rect 72163 35175 72221 35176
rect 72363 35216 72405 35225
rect 72363 35176 72364 35216
rect 72404 35176 72405 35216
rect 72363 35167 72405 35176
rect 72547 35216 72605 35217
rect 72547 35176 72556 35216
rect 72596 35176 72605 35216
rect 72547 35175 72605 35176
rect 74187 35216 74229 35225
rect 74187 35176 74188 35216
rect 74228 35176 74229 35216
rect 74187 35167 74229 35176
rect 74563 35216 74621 35217
rect 74563 35176 74572 35216
rect 74612 35176 74621 35216
rect 74563 35175 74621 35176
rect 75427 35216 75485 35217
rect 75427 35176 75436 35216
rect 75476 35176 75485 35216
rect 75427 35175 75485 35176
rect 77067 35216 77109 35225
rect 77067 35176 77068 35216
rect 77108 35176 77109 35216
rect 77067 35167 77109 35176
rect 77443 35216 77501 35217
rect 77443 35176 77452 35216
rect 77492 35176 77501 35216
rect 77443 35175 77501 35176
rect 78307 35216 78365 35217
rect 78307 35176 78316 35216
rect 78356 35176 78365 35216
rect 78307 35175 78365 35176
rect 55389 35156 55431 35165
rect 51043 35048 51101 35049
rect 51043 35008 51052 35048
rect 51092 35008 51101 35048
rect 51043 35007 51101 35008
rect 52491 35048 52533 35057
rect 52491 35008 52492 35048
rect 52532 35008 52533 35048
rect 52491 34999 52533 35008
rect 58635 35048 58677 35057
rect 58635 35008 58636 35048
rect 58676 35008 58677 35048
rect 58635 34999 58677 35008
rect 63531 35048 63573 35057
rect 63531 35008 63532 35048
rect 63572 35008 63573 35048
rect 63531 34999 63573 35008
rect 64683 35048 64725 35057
rect 64683 35008 64684 35048
rect 64724 35008 64725 35048
rect 64683 34999 64725 35008
rect 67075 35048 67133 35049
rect 67075 35008 67084 35048
rect 67124 35008 67133 35048
rect 67075 35007 67133 35008
rect 71683 35048 71741 35049
rect 71683 35008 71692 35048
rect 71732 35008 71741 35048
rect 71683 35007 71741 35008
rect 72747 35048 72789 35057
rect 72747 35008 72748 35048
rect 72788 35008 72789 35048
rect 72747 34999 72789 35008
rect 46539 34964 46581 34973
rect 46539 34924 46540 34964
rect 46580 34924 46581 34964
rect 46539 34915 46581 34924
rect 48451 34964 48509 34965
rect 48451 34924 48460 34964
rect 48500 34924 48509 34964
rect 48451 34923 48509 34924
rect 52299 34964 52341 34973
rect 52299 34924 52300 34964
rect 52340 34924 52341 34964
rect 52299 34915 52341 34924
rect 57955 34964 58013 34965
rect 57955 34924 57964 34964
rect 58004 34924 58013 34964
rect 57955 34923 58013 34924
rect 58155 34964 58197 34973
rect 58155 34924 58156 34964
rect 58196 34924 58197 34964
rect 58155 34915 58197 34924
rect 62179 34964 62237 34965
rect 62179 34924 62188 34964
rect 62228 34924 62237 34964
rect 62179 34923 62237 34924
rect 62371 34964 62429 34965
rect 62371 34924 62380 34964
rect 62420 34924 62429 34964
rect 62371 34923 62429 34924
rect 69859 34964 69917 34965
rect 69859 34924 69868 34964
rect 69908 34924 69917 34964
rect 69859 34923 69917 34924
rect 71883 34964 71925 34973
rect 71883 34924 71884 34964
rect 71924 34924 71925 34964
rect 71883 34915 71925 34924
rect 72459 34964 72501 34973
rect 72459 34924 72460 34964
rect 72500 34924 72501 34964
rect 72459 34915 72501 34924
rect 76579 34964 76637 34965
rect 76579 34924 76588 34964
rect 76628 34924 76637 34964
rect 76579 34923 76637 34924
rect 79459 34964 79517 34965
rect 79459 34924 79468 34964
rect 79508 34924 79517 34964
rect 79459 34923 79517 34924
rect 576 34796 79584 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 79584 34796
rect 576 34732 79584 34756
rect 50955 34628 50997 34637
rect 50955 34588 50956 34628
rect 50996 34588 50997 34628
rect 50955 34579 50997 34588
rect 55555 34628 55613 34629
rect 55555 34588 55564 34628
rect 55604 34588 55613 34628
rect 55555 34587 55613 34588
rect 66987 34628 67029 34637
rect 66987 34588 66988 34628
rect 67028 34588 67029 34628
rect 66987 34579 67029 34588
rect 68899 34628 68957 34629
rect 68899 34588 68908 34628
rect 68948 34588 68957 34628
rect 68899 34587 68957 34588
rect 77251 34628 77309 34629
rect 77251 34588 77260 34628
rect 77300 34588 77309 34628
rect 77251 34587 77309 34588
rect 45963 34544 46005 34553
rect 45963 34504 45964 34544
rect 46004 34504 46005 34544
rect 45963 34495 46005 34504
rect 49227 34544 49269 34553
rect 49227 34504 49228 34544
rect 49268 34504 49269 34544
rect 49227 34495 49269 34504
rect 51723 34544 51765 34553
rect 51723 34504 51724 34544
rect 51764 34504 51765 34544
rect 51723 34495 51765 34504
rect 52203 34544 52245 34553
rect 52203 34504 52204 34544
rect 52244 34504 52245 34544
rect 52203 34495 52245 34504
rect 52683 34544 52725 34553
rect 52683 34504 52684 34544
rect 52724 34504 52725 34544
rect 52683 34495 52725 34504
rect 56523 34544 56565 34553
rect 56523 34504 56524 34544
rect 56564 34504 56565 34544
rect 56523 34495 56565 34504
rect 57771 34544 57813 34553
rect 57771 34504 57772 34544
rect 57812 34504 57813 34544
rect 57771 34495 57813 34504
rect 61899 34544 61941 34553
rect 61899 34504 61900 34544
rect 61940 34504 61941 34544
rect 61899 34495 61941 34504
rect 66603 34544 66645 34553
rect 66603 34504 66604 34544
rect 66644 34504 66645 34544
rect 66603 34495 66645 34504
rect 67947 34544 67989 34553
rect 67947 34504 67948 34544
rect 67988 34504 67989 34544
rect 67947 34495 67989 34504
rect 71979 34544 72021 34553
rect 71979 34504 71980 34544
rect 72020 34504 72021 34544
rect 71979 34495 72021 34504
rect 77451 34544 77493 34553
rect 77451 34504 77452 34544
rect 77492 34504 77493 34544
rect 77451 34495 77493 34504
rect 78027 34544 78069 34553
rect 78027 34504 78028 34544
rect 78068 34504 78069 34544
rect 78027 34495 78069 34504
rect 46155 34376 46197 34385
rect 46155 34336 46156 34376
rect 46196 34336 46197 34376
rect 46155 34327 46197 34336
rect 46531 34376 46589 34377
rect 46531 34336 46540 34376
rect 46580 34336 46589 34376
rect 46531 34335 46589 34336
rect 47395 34376 47453 34377
rect 47395 34336 47404 34376
rect 47444 34336 47453 34376
rect 47395 34335 47453 34336
rect 49227 34376 49269 34385
rect 49227 34336 49228 34376
rect 49268 34336 49269 34376
rect 49227 34327 49269 34336
rect 49419 34376 49461 34385
rect 49419 34336 49420 34376
rect 49460 34336 49461 34376
rect 49419 34327 49461 34336
rect 49507 34376 49565 34377
rect 49507 34336 49516 34376
rect 49556 34336 49565 34376
rect 49507 34335 49565 34336
rect 50475 34376 50517 34385
rect 50475 34336 50476 34376
rect 50516 34336 50517 34376
rect 50475 34327 50517 34336
rect 50571 34376 50613 34385
rect 50571 34336 50572 34376
rect 50612 34336 50613 34376
rect 50571 34327 50613 34336
rect 50667 34376 50709 34385
rect 50667 34336 50668 34376
rect 50708 34336 50709 34376
rect 50667 34327 50709 34336
rect 50763 34376 50805 34385
rect 50763 34336 50764 34376
rect 50804 34336 50805 34376
rect 50763 34327 50805 34336
rect 50955 34376 50997 34385
rect 50955 34336 50956 34376
rect 50996 34336 50997 34376
rect 50955 34327 50997 34336
rect 51147 34376 51189 34385
rect 51147 34336 51148 34376
rect 51188 34336 51189 34376
rect 51147 34327 51189 34336
rect 51235 34376 51293 34377
rect 51235 34336 51244 34376
rect 51284 34336 51293 34376
rect 51235 34335 51293 34336
rect 51627 34376 51669 34385
rect 51627 34336 51628 34376
rect 51668 34336 51669 34376
rect 51627 34327 51669 34336
rect 51811 34376 51869 34377
rect 51811 34336 51820 34376
rect 51860 34336 51869 34376
rect 51811 34335 51869 34336
rect 52203 34376 52245 34385
rect 52203 34336 52204 34376
rect 52244 34336 52245 34376
rect 52203 34327 52245 34336
rect 52395 34376 52437 34385
rect 52395 34336 52396 34376
rect 52436 34336 52437 34376
rect 52395 34327 52437 34336
rect 52483 34376 52541 34377
rect 52483 34336 52492 34376
rect 52532 34336 52541 34376
rect 52483 34335 52541 34336
rect 53931 34376 53973 34385
rect 53931 34336 53932 34376
rect 53972 34336 53973 34376
rect 53931 34327 53973 34336
rect 54123 34376 54165 34385
rect 54123 34336 54124 34376
rect 54164 34336 54165 34376
rect 54123 34327 54165 34336
rect 54211 34376 54269 34377
rect 54211 34336 54220 34376
rect 54260 34336 54269 34376
rect 54211 34335 54269 34336
rect 54979 34376 55037 34377
rect 54979 34336 54988 34376
rect 55028 34336 55037 34376
rect 54979 34335 55037 34336
rect 55179 34376 55221 34385
rect 55179 34336 55180 34376
rect 55220 34336 55221 34376
rect 55179 34327 55221 34336
rect 55851 34376 55893 34385
rect 55851 34336 55852 34376
rect 55892 34336 55893 34376
rect 55851 34327 55893 34336
rect 55947 34376 55989 34385
rect 55947 34336 55948 34376
rect 55988 34336 55989 34376
rect 55947 34327 55989 34336
rect 56227 34376 56285 34377
rect 56227 34336 56236 34376
rect 56276 34336 56285 34376
rect 56227 34335 56285 34336
rect 57475 34376 57533 34377
rect 57475 34336 57484 34376
rect 57524 34336 57533 34376
rect 57475 34335 57533 34336
rect 57579 34376 57621 34385
rect 57579 34336 57580 34376
rect 57620 34336 57621 34376
rect 57579 34327 57621 34336
rect 57771 34376 57813 34385
rect 57771 34336 57772 34376
rect 57812 34336 57813 34376
rect 57771 34327 57813 34336
rect 57963 34376 58005 34385
rect 57963 34336 57964 34376
rect 58004 34336 58005 34376
rect 57963 34327 58005 34336
rect 58339 34376 58397 34377
rect 58339 34336 58348 34376
rect 58388 34336 58397 34376
rect 58339 34335 58397 34336
rect 59203 34376 59261 34377
rect 59203 34336 59212 34376
rect 59252 34336 59261 34376
rect 59203 34335 59261 34336
rect 61899 34376 61941 34385
rect 61899 34336 61900 34376
rect 61940 34336 61941 34376
rect 61899 34327 61941 34336
rect 62091 34376 62133 34385
rect 62091 34336 62092 34376
rect 62132 34336 62133 34376
rect 62091 34327 62133 34336
rect 62179 34376 62237 34377
rect 62179 34336 62188 34376
rect 62228 34336 62237 34376
rect 62179 34335 62237 34336
rect 62571 34376 62613 34385
rect 62571 34336 62572 34376
rect 62612 34336 62613 34376
rect 62571 34327 62613 34336
rect 62763 34376 62805 34385
rect 62763 34336 62764 34376
rect 62804 34336 62805 34376
rect 62763 34327 62805 34336
rect 62851 34376 62909 34377
rect 62851 34336 62860 34376
rect 62900 34336 62909 34376
rect 62851 34335 62909 34336
rect 63427 34376 63485 34377
rect 63427 34336 63436 34376
rect 63476 34336 63485 34376
rect 63427 34335 63485 34336
rect 64291 34376 64349 34377
rect 64291 34336 64300 34376
rect 64340 34336 64349 34376
rect 64291 34335 64349 34336
rect 66123 34376 66165 34385
rect 66123 34336 66124 34376
rect 66164 34336 66165 34376
rect 66123 34327 66165 34336
rect 66315 34376 66357 34385
rect 66315 34336 66316 34376
rect 66356 34336 66357 34376
rect 66315 34327 66357 34336
rect 66403 34376 66461 34377
rect 66403 34336 66412 34376
rect 66452 34336 66461 34376
rect 66403 34335 66461 34336
rect 66987 34376 67029 34385
rect 66987 34336 66988 34376
rect 67028 34336 67029 34376
rect 66987 34327 67029 34336
rect 67179 34376 67221 34385
rect 67179 34336 67180 34376
rect 67220 34336 67221 34376
rect 67179 34327 67221 34336
rect 67267 34376 67325 34377
rect 67267 34336 67276 34376
rect 67316 34336 67325 34376
rect 67267 34335 67325 34336
rect 67459 34376 67517 34377
rect 67459 34336 67468 34376
rect 67508 34336 67517 34376
rect 67459 34335 67517 34336
rect 67563 34376 67605 34385
rect 67563 34336 67564 34376
rect 67604 34336 67605 34376
rect 67563 34327 67605 34336
rect 67668 34376 67710 34385
rect 67668 34336 67669 34376
rect 67709 34336 67710 34376
rect 67668 34327 67710 34336
rect 70051 34376 70109 34377
rect 70051 34336 70060 34376
rect 70100 34336 70109 34376
rect 70051 34335 70109 34336
rect 70915 34376 70973 34377
rect 70915 34336 70924 34376
rect 70964 34336 70973 34376
rect 70915 34335 70973 34336
rect 71307 34376 71349 34385
rect 71307 34336 71308 34376
rect 71348 34336 71349 34376
rect 71307 34327 71349 34336
rect 71683 34376 71741 34377
rect 71683 34336 71692 34376
rect 71732 34336 71741 34376
rect 71683 34335 71741 34336
rect 71787 34376 71829 34385
rect 71787 34336 71788 34376
rect 71828 34336 71829 34376
rect 71787 34327 71829 34336
rect 71979 34376 72021 34385
rect 71979 34336 71980 34376
rect 72020 34336 72021 34376
rect 71979 34327 72021 34336
rect 72171 34376 72213 34385
rect 72171 34336 72172 34376
rect 72212 34336 72213 34376
rect 72171 34327 72213 34336
rect 72547 34376 72605 34377
rect 72547 34336 72556 34376
rect 72596 34336 72605 34376
rect 72547 34335 72605 34336
rect 73452 34376 73494 34385
rect 73452 34336 73453 34376
rect 73493 34336 73494 34376
rect 73452 34327 73494 34336
rect 76011 34376 76053 34385
rect 76011 34336 76012 34376
rect 76052 34336 76053 34376
rect 76011 34327 76053 34336
rect 76203 34376 76245 34385
rect 76203 34336 76204 34376
rect 76244 34336 76245 34376
rect 76203 34327 76245 34336
rect 76291 34376 76349 34377
rect 76291 34336 76300 34376
rect 76340 34336 76349 34376
rect 76291 34335 76349 34336
rect 76579 34376 76637 34377
rect 76579 34336 76588 34376
rect 76628 34336 76637 34376
rect 76579 34335 76637 34336
rect 76875 34376 76917 34385
rect 76875 34336 76876 34376
rect 76916 34336 76917 34376
rect 76875 34327 76917 34336
rect 76971 34376 77013 34385
rect 76971 34336 76972 34376
rect 77012 34336 77013 34376
rect 76971 34327 77013 34336
rect 77451 34376 77493 34385
rect 77451 34336 77452 34376
rect 77492 34336 77493 34376
rect 77451 34327 77493 34336
rect 77643 34376 77685 34385
rect 77643 34336 77644 34376
rect 77684 34336 77685 34376
rect 77643 34327 77685 34336
rect 77731 34376 77789 34377
rect 77731 34336 77740 34376
rect 77780 34336 77789 34376
rect 77731 34335 77789 34336
rect 77923 34376 77981 34377
rect 77923 34336 77932 34376
rect 77972 34336 77981 34376
rect 77923 34335 77981 34336
rect 78123 34376 78165 34385
rect 78123 34336 78124 34376
rect 78164 34336 78165 34376
rect 78123 34327 78165 34336
rect 55083 34292 55125 34301
rect 55083 34252 55084 34292
rect 55124 34252 55125 34292
rect 55083 34243 55125 34252
rect 62667 34292 62709 34301
rect 62667 34252 62668 34292
rect 62708 34252 62709 34292
rect 62667 34243 62709 34252
rect 63051 34292 63093 34301
rect 63051 34252 63052 34292
rect 63092 34252 63093 34292
rect 63051 34243 63093 34252
rect 76107 34292 76149 34301
rect 76107 34252 76108 34292
rect 76148 34252 76149 34292
rect 76107 34243 76149 34252
rect 48547 34208 48605 34209
rect 48547 34168 48556 34208
rect 48596 34168 48605 34208
rect 48547 34167 48605 34168
rect 54019 34208 54077 34209
rect 54019 34168 54028 34208
rect 54068 34168 54077 34208
rect 54019 34167 54077 34168
rect 60355 34208 60413 34209
rect 60355 34168 60364 34208
rect 60404 34168 60413 34208
rect 60355 34167 60413 34168
rect 65443 34208 65501 34209
rect 65443 34168 65452 34208
rect 65492 34168 65501 34208
rect 65443 34167 65501 34168
rect 66211 34208 66269 34209
rect 66211 34168 66220 34208
rect 66260 34168 66269 34208
rect 66211 34167 66269 34168
rect 74563 34208 74621 34209
rect 74563 34168 74572 34208
rect 74612 34168 74621 34208
rect 74563 34167 74621 34168
rect 576 34040 79584 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 79584 34040
rect 576 33976 79584 34000
rect 46435 33872 46493 33873
rect 46435 33832 46444 33872
rect 46484 33832 46493 33872
rect 46435 33831 46493 33832
rect 58339 33872 58397 33873
rect 58339 33832 58348 33872
rect 58388 33832 58397 33872
rect 58339 33831 58397 33832
rect 76771 33872 76829 33873
rect 76771 33832 76780 33872
rect 76820 33832 76829 33872
rect 76771 33831 76829 33832
rect 52203 33788 52245 33797
rect 52203 33748 52204 33788
rect 52244 33748 52245 33788
rect 52203 33739 52245 33748
rect 55275 33788 55317 33797
rect 55275 33748 55276 33788
rect 55316 33748 55317 33788
rect 55275 33739 55317 33748
rect 62283 33788 62325 33797
rect 62283 33748 62284 33788
rect 62324 33748 62325 33788
rect 62283 33739 62325 33748
rect 62763 33788 62805 33797
rect 62763 33748 62764 33788
rect 62804 33748 62805 33788
rect 62763 33739 62805 33748
rect 63147 33788 63189 33797
rect 63147 33748 63148 33788
rect 63188 33748 63189 33788
rect 63147 33739 63189 33748
rect 71691 33788 71733 33797
rect 71691 33748 71692 33788
rect 71732 33748 71733 33788
rect 71691 33739 71733 33748
rect 46539 33704 46581 33713
rect 46539 33664 46540 33704
rect 46580 33664 46581 33704
rect 46539 33655 46581 33664
rect 46635 33704 46677 33713
rect 46635 33664 46636 33704
rect 46676 33664 46677 33704
rect 46635 33655 46677 33664
rect 46731 33704 46773 33713
rect 46731 33664 46732 33704
rect 46772 33664 46773 33704
rect 46731 33655 46773 33664
rect 48939 33704 48981 33713
rect 48939 33664 48940 33704
rect 48980 33664 48981 33704
rect 48939 33655 48981 33664
rect 49131 33704 49173 33713
rect 49131 33664 49132 33704
rect 49172 33664 49173 33704
rect 49131 33655 49173 33664
rect 49219 33704 49277 33705
rect 49219 33664 49228 33704
rect 49268 33664 49277 33704
rect 49219 33663 49277 33664
rect 52579 33704 52637 33705
rect 52579 33664 52588 33704
rect 52628 33664 52637 33704
rect 52579 33663 52637 33664
rect 53443 33704 53501 33705
rect 53443 33664 53452 33704
rect 53492 33664 53501 33704
rect 53443 33663 53501 33664
rect 54883 33704 54941 33705
rect 54883 33664 54892 33704
rect 54932 33664 54941 33704
rect 54883 33663 54941 33664
rect 55179 33704 55221 33713
rect 55179 33664 55180 33704
rect 55220 33664 55221 33704
rect 55179 33655 55221 33664
rect 58443 33704 58485 33713
rect 58443 33664 58444 33704
rect 58484 33664 58485 33704
rect 58443 33655 58485 33664
rect 58539 33704 58581 33713
rect 58539 33664 58540 33704
rect 58580 33664 58581 33704
rect 58819 33704 58877 33705
rect 58539 33655 58581 33664
rect 58635 33659 58677 33668
rect 58819 33664 58828 33704
rect 58868 33664 58877 33704
rect 58819 33663 58877 33664
rect 59019 33704 59061 33713
rect 59019 33664 59020 33704
rect 59060 33664 59061 33704
rect 54603 33620 54645 33629
rect 54603 33580 54604 33620
rect 54644 33580 54645 33620
rect 58635 33619 58636 33659
rect 58676 33619 58677 33659
rect 59019 33655 59061 33664
rect 62187 33704 62229 33713
rect 62187 33664 62188 33704
rect 62228 33664 62229 33704
rect 62187 33655 62229 33664
rect 62379 33704 62421 33713
rect 62379 33664 62380 33704
rect 62420 33664 62421 33704
rect 62379 33655 62421 33664
rect 62467 33704 62525 33705
rect 62467 33664 62476 33704
rect 62516 33664 62525 33704
rect 62467 33663 62525 33664
rect 62667 33704 62709 33713
rect 62667 33664 62668 33704
rect 62708 33664 62709 33704
rect 62667 33655 62709 33664
rect 62851 33704 62909 33705
rect 62851 33664 62860 33704
rect 62900 33664 62909 33704
rect 62851 33663 62909 33664
rect 63043 33704 63101 33705
rect 63043 33664 63052 33704
rect 63092 33664 63101 33704
rect 63043 33663 63101 33664
rect 63243 33704 63285 33713
rect 63243 33664 63244 33704
rect 63284 33664 63285 33704
rect 63243 33655 63285 33664
rect 66219 33704 66261 33713
rect 66219 33664 66220 33704
rect 66260 33664 66261 33704
rect 66219 33655 66261 33664
rect 66595 33704 66653 33705
rect 66595 33664 66604 33704
rect 66644 33664 66653 33704
rect 66595 33663 66653 33664
rect 67459 33704 67517 33705
rect 67459 33664 67468 33704
rect 67508 33664 67517 33704
rect 67459 33663 67517 33664
rect 71587 33704 71645 33705
rect 71587 33664 71596 33704
rect 71636 33664 71645 33704
rect 71587 33663 71645 33664
rect 71787 33704 71829 33713
rect 71787 33664 71788 33704
rect 71828 33664 71829 33704
rect 71787 33655 71829 33664
rect 71979 33704 72021 33713
rect 71979 33664 71980 33704
rect 72020 33664 72021 33704
rect 71979 33655 72021 33664
rect 72171 33704 72213 33713
rect 72171 33664 72172 33704
rect 72212 33664 72213 33704
rect 72171 33655 72213 33664
rect 72259 33704 72317 33705
rect 72259 33664 72268 33704
rect 72308 33664 72317 33704
rect 72259 33663 72317 33664
rect 72451 33704 72509 33705
rect 72451 33664 72460 33704
rect 72500 33664 72509 33704
rect 72451 33663 72509 33664
rect 72651 33704 72693 33713
rect 72651 33664 72652 33704
rect 72692 33664 72693 33704
rect 72651 33655 72693 33664
rect 75715 33704 75773 33705
rect 75715 33664 75724 33704
rect 75764 33664 75773 33704
rect 75715 33663 75773 33664
rect 75819 33704 75861 33713
rect 75819 33664 75820 33704
rect 75860 33664 75861 33704
rect 75819 33655 75861 33664
rect 76011 33704 76053 33713
rect 76011 33664 76012 33704
rect 76052 33664 76053 33704
rect 76011 33655 76053 33664
rect 76203 33704 76245 33713
rect 76203 33664 76204 33704
rect 76244 33664 76245 33704
rect 76203 33655 76245 33664
rect 76299 33704 76341 33713
rect 76299 33664 76300 33704
rect 76340 33664 76341 33704
rect 76299 33655 76341 33664
rect 76395 33704 76437 33713
rect 76395 33664 76396 33704
rect 76436 33664 76437 33704
rect 76395 33655 76437 33664
rect 76491 33704 76533 33713
rect 76491 33664 76492 33704
rect 76532 33664 76533 33704
rect 76491 33655 76533 33664
rect 76683 33704 76725 33713
rect 76683 33664 76684 33704
rect 76724 33664 76725 33704
rect 76683 33655 76725 33664
rect 76875 33704 76917 33713
rect 76875 33664 76876 33704
rect 76916 33664 76917 33704
rect 76875 33655 76917 33664
rect 76963 33704 77021 33705
rect 76963 33664 76972 33704
rect 77012 33664 77021 33704
rect 76963 33663 77021 33664
rect 77259 33704 77301 33713
rect 77259 33664 77260 33704
rect 77300 33664 77301 33704
rect 77259 33655 77301 33664
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77451 33655 77493 33664
rect 77539 33704 77597 33705
rect 77539 33664 77548 33704
rect 77588 33664 77597 33704
rect 77539 33663 77597 33664
rect 58635 33610 58677 33619
rect 72555 33620 72597 33629
rect 54603 33571 54645 33580
rect 72555 33580 72556 33620
rect 72596 33580 72597 33620
rect 72555 33571 72597 33580
rect 46251 33536 46293 33545
rect 46251 33496 46252 33536
rect 46292 33496 46293 33536
rect 46251 33487 46293 33496
rect 55555 33536 55613 33537
rect 55555 33496 55564 33536
rect 55604 33496 55613 33536
rect 55555 33495 55613 33496
rect 56139 33536 56181 33545
rect 56139 33496 56140 33536
rect 56180 33496 56181 33536
rect 56139 33487 56181 33496
rect 59211 33536 59253 33545
rect 59211 33496 59212 33536
rect 59252 33496 59253 33536
rect 59211 33487 59253 33496
rect 63723 33536 63765 33545
rect 63723 33496 63724 33536
rect 63764 33496 63765 33536
rect 63723 33487 63765 33496
rect 69771 33536 69813 33545
rect 69771 33496 69772 33536
rect 69812 33496 69813 33536
rect 69771 33487 69813 33496
rect 75051 33536 75093 33545
rect 75051 33496 75052 33536
rect 75092 33496 75093 33536
rect 75051 33487 75093 33496
rect 77835 33536 77877 33545
rect 77835 33496 77836 33536
rect 77876 33496 77877 33536
rect 77835 33487 77877 33496
rect 48939 33452 48981 33461
rect 48939 33412 48940 33452
rect 48980 33412 48981 33452
rect 48939 33403 48981 33412
rect 58923 33452 58965 33461
rect 58923 33412 58924 33452
rect 58964 33412 58965 33452
rect 58923 33403 58965 33412
rect 68611 33452 68669 33453
rect 68611 33412 68620 33452
rect 68660 33412 68669 33452
rect 68611 33411 68669 33412
rect 71979 33452 72021 33461
rect 71979 33412 71980 33452
rect 72020 33412 72021 33452
rect 71979 33403 72021 33412
rect 76011 33452 76053 33461
rect 76011 33412 76012 33452
rect 76052 33412 76053 33452
rect 76011 33403 76053 33412
rect 77259 33452 77301 33461
rect 77259 33412 77260 33452
rect 77300 33412 77301 33452
rect 77259 33403 77301 33412
rect 576 33284 79584 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 75112 33284
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75480 33244 79584 33284
rect 576 33220 79584 33244
rect 42987 33116 43029 33125
rect 42987 33076 42988 33116
rect 43028 33076 43029 33116
rect 42987 33067 43029 33076
rect 47595 33116 47637 33125
rect 47595 33076 47596 33116
rect 47636 33076 47637 33116
rect 47595 33067 47637 33076
rect 66507 33116 66549 33125
rect 66507 33076 66508 33116
rect 66548 33076 66549 33116
rect 66507 33067 66549 33076
rect 77155 33116 77213 33117
rect 77155 33076 77164 33116
rect 77204 33076 77213 33116
rect 77155 33075 77213 33076
rect 43947 33032 43989 33041
rect 43947 32992 43948 33032
rect 43988 32992 43989 33032
rect 43947 32983 43989 32992
rect 46915 33032 46973 33033
rect 46915 32992 46924 33032
rect 46964 32992 46973 33032
rect 46915 32991 46973 32992
rect 48075 33032 48117 33041
rect 48075 32992 48076 33032
rect 48116 32992 48117 33032
rect 48075 32983 48117 32992
rect 51627 33032 51669 33041
rect 51627 32992 51628 33032
rect 51668 32992 51669 33032
rect 51627 32983 51669 32992
rect 55467 33032 55509 33041
rect 55467 32992 55468 33032
rect 55508 32992 55509 33032
rect 55467 32983 55509 32992
rect 61323 33032 61365 33041
rect 61323 32992 61324 33032
rect 61364 32992 61365 33032
rect 61323 32983 61365 32992
rect 78115 33032 78173 33033
rect 78115 32992 78124 33032
rect 78164 32992 78173 33032
rect 78115 32991 78173 32992
rect 78411 33032 78453 33041
rect 78411 32992 78412 33032
rect 78452 32992 78453 33032
rect 78411 32983 78453 32992
rect 42787 32948 42845 32949
rect 42787 32908 42796 32948
rect 42836 32908 42845 32948
rect 42787 32907 42845 32908
rect 45675 32864 45717 32873
rect 45675 32824 45676 32864
rect 45716 32824 45717 32864
rect 45675 32815 45717 32824
rect 45867 32864 45909 32873
rect 45867 32824 45868 32864
rect 45908 32824 45909 32864
rect 45867 32815 45909 32824
rect 45955 32864 46013 32865
rect 45955 32824 45964 32864
rect 46004 32824 46013 32864
rect 45955 32823 46013 32824
rect 46243 32864 46301 32865
rect 46243 32824 46252 32864
rect 46292 32824 46301 32864
rect 46243 32823 46301 32824
rect 46539 32864 46581 32873
rect 46539 32824 46540 32864
rect 46580 32824 46581 32864
rect 46539 32815 46581 32824
rect 46635 32864 46677 32873
rect 46635 32824 46636 32864
rect 46676 32824 46677 32864
rect 46635 32815 46677 32824
rect 47107 32864 47165 32865
rect 47107 32824 47116 32864
rect 47156 32824 47165 32864
rect 47107 32823 47165 32824
rect 47307 32864 47349 32873
rect 47307 32824 47308 32864
rect 47348 32824 47349 32864
rect 47307 32815 47349 32824
rect 47491 32864 47549 32865
rect 47491 32824 47500 32864
rect 47540 32824 47549 32864
rect 47491 32823 47549 32824
rect 47691 32864 47733 32873
rect 47691 32824 47692 32864
rect 47732 32824 47733 32864
rect 47691 32815 47733 32824
rect 48267 32864 48309 32873
rect 48267 32824 48268 32864
rect 48308 32824 48309 32864
rect 48267 32815 48309 32824
rect 48643 32864 48701 32865
rect 48643 32824 48652 32864
rect 48692 32824 48701 32864
rect 48643 32823 48701 32824
rect 49507 32864 49565 32865
rect 49507 32824 49516 32864
rect 49556 32824 49565 32864
rect 49507 32823 49565 32824
rect 50851 32864 50909 32865
rect 50851 32824 50860 32864
rect 50900 32824 50909 32864
rect 50851 32823 50909 32824
rect 51051 32864 51093 32873
rect 51051 32824 51052 32864
rect 51092 32824 51093 32864
rect 51051 32815 51093 32824
rect 51243 32864 51285 32873
rect 51243 32824 51244 32864
rect 51284 32824 51285 32864
rect 51243 32815 51285 32824
rect 51427 32864 51485 32865
rect 51427 32824 51436 32864
rect 51476 32824 51485 32864
rect 51427 32823 51485 32824
rect 53643 32864 53685 32873
rect 53643 32824 53644 32864
rect 53684 32824 53685 32864
rect 53643 32815 53685 32824
rect 53739 32864 53781 32873
rect 53739 32824 53740 32864
rect 53780 32824 53781 32864
rect 53739 32815 53781 32824
rect 53835 32864 53877 32873
rect 53835 32824 53836 32864
rect 53876 32824 53877 32864
rect 53835 32815 53877 32824
rect 53931 32864 53973 32873
rect 53931 32824 53932 32864
rect 53972 32824 53973 32864
rect 53931 32815 53973 32824
rect 54787 32864 54845 32865
rect 54787 32824 54796 32864
rect 54836 32824 54845 32864
rect 54787 32823 54845 32824
rect 54891 32864 54933 32873
rect 54891 32824 54892 32864
rect 54932 32824 54933 32864
rect 54891 32815 54933 32824
rect 54987 32864 55029 32873
rect 54987 32824 54988 32864
rect 55028 32824 55029 32864
rect 54987 32815 55029 32824
rect 55171 32864 55229 32865
rect 55171 32824 55180 32864
rect 55220 32824 55229 32864
rect 55171 32823 55229 32824
rect 55275 32864 55317 32873
rect 55275 32824 55276 32864
rect 55316 32824 55317 32864
rect 55275 32815 55317 32824
rect 55467 32864 55509 32873
rect 55467 32824 55468 32864
rect 55508 32824 55509 32864
rect 55467 32815 55509 32824
rect 55659 32864 55701 32873
rect 55659 32824 55660 32864
rect 55700 32824 55701 32864
rect 55659 32815 55701 32824
rect 56035 32864 56093 32865
rect 56035 32824 56044 32864
rect 56084 32824 56093 32864
rect 56035 32823 56093 32824
rect 56899 32864 56957 32865
rect 56899 32824 56908 32864
rect 56948 32824 56957 32864
rect 56899 32823 56957 32824
rect 58251 32864 58293 32873
rect 58251 32824 58252 32864
rect 58292 32824 58293 32864
rect 58251 32815 58293 32824
rect 58443 32864 58485 32873
rect 58443 32824 58444 32864
rect 58484 32824 58485 32864
rect 58443 32815 58485 32824
rect 58531 32864 58589 32865
rect 58531 32824 58540 32864
rect 58580 32824 58589 32864
rect 58531 32823 58589 32824
rect 59107 32864 59165 32865
rect 59107 32824 59116 32864
rect 59156 32824 59165 32864
rect 59107 32823 59165 32824
rect 59971 32864 60029 32865
rect 59971 32824 59980 32864
rect 60020 32824 60029 32864
rect 59971 32823 60029 32824
rect 62475 32864 62517 32873
rect 62475 32824 62476 32864
rect 62516 32824 62517 32864
rect 62475 32815 62517 32824
rect 62571 32864 62613 32873
rect 62571 32824 62572 32864
rect 62612 32824 62613 32864
rect 62571 32815 62613 32824
rect 62667 32864 62709 32873
rect 62667 32824 62668 32864
rect 62708 32824 62709 32864
rect 62667 32815 62709 32824
rect 63619 32864 63677 32865
rect 63619 32824 63628 32864
rect 63668 32824 63677 32864
rect 63619 32823 63677 32824
rect 64483 32864 64541 32865
rect 64483 32824 64492 32864
rect 64532 32824 64541 32864
rect 64483 32823 64541 32824
rect 66027 32864 66069 32873
rect 66027 32824 66028 32864
rect 66068 32824 66069 32864
rect 66027 32815 66069 32824
rect 66123 32864 66165 32873
rect 66123 32824 66124 32864
rect 66164 32824 66165 32864
rect 66123 32815 66165 32824
rect 66219 32864 66261 32873
rect 66219 32824 66220 32864
rect 66260 32824 66261 32864
rect 66219 32815 66261 32824
rect 66315 32864 66357 32873
rect 66315 32824 66316 32864
rect 66356 32824 66357 32864
rect 66315 32815 66357 32824
rect 66507 32864 66549 32873
rect 66507 32824 66508 32864
rect 66548 32824 66549 32864
rect 66507 32815 66549 32824
rect 66699 32864 66741 32873
rect 66699 32824 66700 32864
rect 66740 32824 66741 32864
rect 66699 32815 66741 32824
rect 66787 32864 66845 32865
rect 66787 32824 66796 32864
rect 66836 32824 66845 32864
rect 66787 32823 66845 32824
rect 68803 32864 68861 32865
rect 68803 32824 68812 32864
rect 68852 32824 68861 32864
rect 68803 32823 68861 32824
rect 68907 32864 68949 32873
rect 68907 32824 68908 32864
rect 68948 32824 68949 32864
rect 68907 32815 68949 32824
rect 69099 32864 69141 32873
rect 69099 32824 69100 32864
rect 69140 32824 69141 32864
rect 69099 32815 69141 32824
rect 69667 32864 69725 32865
rect 69667 32824 69676 32864
rect 69716 32824 69725 32864
rect 69667 32823 69725 32824
rect 70531 32864 70589 32865
rect 70531 32824 70540 32864
rect 70580 32824 70589 32864
rect 70531 32823 70589 32824
rect 72171 32864 72213 32873
rect 72171 32824 72172 32864
rect 72212 32824 72213 32864
rect 72171 32815 72213 32824
rect 72547 32864 72605 32865
rect 72547 32824 72556 32864
rect 72596 32824 72605 32864
rect 74763 32864 74805 32873
rect 72547 32823 72605 32824
rect 73411 32853 73469 32854
rect 73411 32813 73420 32853
rect 73460 32813 73469 32853
rect 74763 32824 74764 32864
rect 74804 32824 74805 32864
rect 74763 32815 74805 32824
rect 75139 32864 75197 32865
rect 75139 32824 75148 32864
rect 75188 32824 75197 32864
rect 75139 32823 75197 32824
rect 76003 32864 76061 32865
rect 76003 32824 76012 32864
rect 76052 32824 76061 32864
rect 76003 32823 76061 32824
rect 77443 32864 77501 32865
rect 77443 32824 77452 32864
rect 77492 32824 77501 32864
rect 77443 32823 77501 32824
rect 77739 32864 77781 32873
rect 77739 32824 77740 32864
rect 77780 32824 77781 32864
rect 77739 32815 77781 32824
rect 77835 32864 77877 32873
rect 77835 32824 77836 32864
rect 77876 32824 77877 32864
rect 77835 32815 77877 32824
rect 78307 32864 78365 32865
rect 78307 32824 78316 32864
rect 78356 32824 78365 32864
rect 78307 32823 78365 32824
rect 78507 32864 78549 32873
rect 78507 32824 78508 32864
rect 78548 32824 78549 32864
rect 78507 32815 78549 32824
rect 73411 32812 73469 32813
rect 47211 32780 47253 32789
rect 47211 32740 47212 32780
rect 47252 32740 47253 32780
rect 47211 32731 47253 32740
rect 50955 32780 50997 32789
rect 50955 32740 50956 32780
rect 50996 32740 50997 32780
rect 50955 32731 50997 32740
rect 51339 32780 51381 32789
rect 51339 32740 51340 32780
rect 51380 32740 51381 32780
rect 51339 32731 51381 32740
rect 58347 32780 58389 32789
rect 58347 32740 58348 32780
rect 58388 32740 58389 32780
rect 58347 32731 58389 32740
rect 58731 32780 58773 32789
rect 58731 32740 58732 32780
rect 58772 32740 58773 32780
rect 58731 32731 58773 32740
rect 63243 32780 63285 32789
rect 63243 32740 63244 32780
rect 63284 32740 63285 32780
rect 63243 32731 63285 32740
rect 69291 32780 69333 32789
rect 69291 32740 69292 32780
rect 69332 32740 69333 32780
rect 69291 32731 69333 32740
rect 45763 32696 45821 32697
rect 45763 32656 45772 32696
rect 45812 32656 45821 32696
rect 45763 32655 45821 32656
rect 50659 32696 50717 32697
rect 50659 32656 50668 32696
rect 50708 32656 50717 32696
rect 50659 32655 50717 32656
rect 58051 32696 58109 32697
rect 58051 32656 58060 32696
rect 58100 32656 58109 32696
rect 58051 32655 58109 32656
rect 61123 32696 61181 32697
rect 61123 32656 61132 32696
rect 61172 32656 61181 32696
rect 61123 32655 61181 32656
rect 62371 32696 62429 32697
rect 62371 32656 62380 32696
rect 62420 32656 62429 32696
rect 62371 32655 62429 32656
rect 65635 32696 65693 32697
rect 65635 32656 65644 32696
rect 65684 32656 65693 32696
rect 65635 32655 65693 32656
rect 68995 32696 69053 32697
rect 68995 32656 69004 32696
rect 69044 32656 69053 32696
rect 68995 32655 69053 32656
rect 71683 32696 71741 32697
rect 71683 32656 71692 32696
rect 71732 32656 71741 32696
rect 71683 32655 71741 32656
rect 74563 32696 74621 32697
rect 74563 32656 74572 32696
rect 74612 32656 74621 32696
rect 74563 32655 74621 32656
rect 576 32528 79584 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 76352 32528
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76720 32488 79584 32528
rect 576 32464 79584 32488
rect 48259 32360 48317 32361
rect 48259 32320 48268 32360
rect 48308 32320 48317 32360
rect 48259 32319 48317 32320
rect 48739 32360 48797 32361
rect 48739 32320 48748 32360
rect 48788 32320 48797 32360
rect 48739 32319 48797 32320
rect 54211 32360 54269 32361
rect 54211 32320 54220 32360
rect 54260 32320 54269 32360
rect 54211 32319 54269 32320
rect 62755 32360 62813 32361
rect 62755 32320 62764 32360
rect 62804 32320 62813 32360
rect 62755 32319 62813 32320
rect 69955 32360 70013 32361
rect 69955 32320 69964 32360
rect 70004 32320 70013 32360
rect 69955 32319 70013 32320
rect 75907 32360 75965 32361
rect 75907 32320 75916 32360
rect 75956 32320 75965 32360
rect 75907 32319 75965 32320
rect 45867 32276 45909 32285
rect 45867 32236 45868 32276
rect 45908 32236 45909 32276
rect 45867 32227 45909 32236
rect 58731 32276 58773 32285
rect 58731 32236 58732 32276
rect 58772 32236 58773 32276
rect 58731 32227 58773 32236
rect 63435 32276 63477 32285
rect 63435 32236 63436 32276
rect 63476 32236 63477 32276
rect 63339 32219 63381 32228
rect 63435 32227 63477 32236
rect 66027 32276 66069 32285
rect 66027 32236 66028 32276
rect 66068 32236 66069 32276
rect 66027 32227 66069 32236
rect 71979 32276 72021 32285
rect 71979 32236 71980 32276
rect 72020 32236 72021 32276
rect 71979 32227 72021 32236
rect 76779 32276 76821 32285
rect 76779 32236 76780 32276
rect 76820 32236 76821 32276
rect 76779 32227 76821 32236
rect 77067 32276 77109 32285
rect 77067 32236 77068 32276
rect 77108 32236 77109 32276
rect 77067 32227 77109 32236
rect 42411 32192 42453 32201
rect 42411 32152 42412 32192
rect 42452 32152 42453 32192
rect 42411 32143 42453 32152
rect 42507 32192 42549 32201
rect 42507 32152 42508 32192
rect 42548 32152 42549 32192
rect 42507 32143 42549 32152
rect 42603 32192 42645 32201
rect 42603 32152 42604 32192
rect 42644 32152 42645 32192
rect 42603 32143 42645 32152
rect 42699 32192 42741 32201
rect 42699 32152 42700 32192
rect 42740 32152 42741 32192
rect 42699 32143 42741 32152
rect 42891 32192 42933 32201
rect 42891 32152 42892 32192
rect 42932 32152 42933 32192
rect 42891 32143 42933 32152
rect 43075 32192 43133 32193
rect 43075 32152 43084 32192
rect 43124 32152 43133 32192
rect 43075 32151 43133 32152
rect 43275 32192 43317 32201
rect 43275 32152 43276 32192
rect 43316 32152 43317 32192
rect 43275 32143 43317 32152
rect 43651 32192 43709 32193
rect 43651 32152 43660 32192
rect 43700 32152 43709 32192
rect 43651 32151 43709 32152
rect 44515 32192 44573 32193
rect 44515 32152 44524 32192
rect 44564 32152 44573 32192
rect 44515 32151 44573 32152
rect 46243 32192 46301 32193
rect 46243 32152 46252 32192
rect 46292 32152 46301 32192
rect 46243 32151 46301 32152
rect 47107 32192 47165 32193
rect 47107 32152 47116 32192
rect 47156 32152 47165 32192
rect 47107 32151 47165 32152
rect 48451 32192 48509 32193
rect 48451 32152 48460 32192
rect 48500 32152 48509 32192
rect 48451 32151 48509 32152
rect 48843 32192 48885 32201
rect 48843 32152 48844 32192
rect 48884 32152 48885 32192
rect 48843 32143 48885 32152
rect 48939 32192 48981 32201
rect 48939 32152 48940 32192
rect 48980 32152 48981 32192
rect 49419 32192 49461 32201
rect 48939 32143 48981 32152
rect 49035 32147 49077 32156
rect 49035 32107 49036 32147
rect 49076 32107 49077 32147
rect 49419 32152 49420 32192
rect 49460 32152 49461 32192
rect 49419 32143 49461 32152
rect 51147 32192 51189 32201
rect 51147 32152 51148 32192
rect 51188 32152 51189 32192
rect 51147 32143 51189 32152
rect 51523 32192 51581 32193
rect 51523 32152 51532 32192
rect 51572 32152 51581 32192
rect 51523 32151 51581 32152
rect 52387 32192 52445 32193
rect 52387 32152 52396 32192
rect 52436 32152 52445 32192
rect 52387 32151 52445 32152
rect 54123 32192 54165 32201
rect 54123 32152 54124 32192
rect 54164 32152 54165 32192
rect 54123 32143 54165 32152
rect 54315 32192 54357 32201
rect 54315 32152 54316 32192
rect 54356 32152 54357 32192
rect 54315 32143 54357 32152
rect 54403 32192 54461 32193
rect 54403 32152 54412 32192
rect 54452 32152 54461 32192
rect 54403 32151 54461 32152
rect 54603 32192 54645 32201
rect 54603 32152 54604 32192
rect 54644 32152 54645 32192
rect 54603 32143 54645 32152
rect 54699 32192 54741 32201
rect 54699 32152 54700 32192
rect 54740 32152 54741 32192
rect 54699 32143 54741 32152
rect 54795 32192 54837 32201
rect 54795 32152 54796 32192
rect 54836 32152 54837 32192
rect 54795 32143 54837 32152
rect 54891 32192 54933 32201
rect 54891 32152 54892 32192
rect 54932 32152 54933 32192
rect 54891 32143 54933 32152
rect 58339 32192 58397 32193
rect 58339 32152 58348 32192
rect 58388 32152 58397 32192
rect 58339 32151 58397 32152
rect 58635 32192 58677 32201
rect 58635 32152 58636 32192
rect 58676 32152 58677 32192
rect 58635 32143 58677 32152
rect 59211 32192 59253 32201
rect 59211 32152 59212 32192
rect 59252 32152 59253 32192
rect 59211 32143 59253 32152
rect 59395 32192 59453 32193
rect 59395 32152 59404 32192
rect 59444 32152 59453 32192
rect 59395 32151 59453 32152
rect 59587 32192 59645 32193
rect 59587 32152 59596 32192
rect 59636 32152 59645 32192
rect 59587 32151 59645 32152
rect 59691 32192 59733 32201
rect 59691 32152 59692 32192
rect 59732 32152 59733 32192
rect 59691 32143 59733 32152
rect 59883 32192 59925 32201
rect 59883 32152 59884 32192
rect 59924 32152 59925 32192
rect 59883 32143 59925 32152
rect 60363 32192 60405 32201
rect 60363 32152 60364 32192
rect 60404 32152 60405 32192
rect 60363 32143 60405 32152
rect 60739 32192 60797 32193
rect 60739 32152 60748 32192
rect 60788 32152 60797 32192
rect 60739 32151 60797 32152
rect 61603 32192 61661 32193
rect 61603 32152 61612 32192
rect 61652 32152 61661 32192
rect 61603 32151 61661 32152
rect 63043 32192 63101 32193
rect 63043 32152 63052 32192
rect 63092 32152 63101 32192
rect 63339 32179 63340 32219
rect 63380 32179 63381 32219
rect 64099 32213 64157 32214
rect 63339 32170 63381 32179
rect 63915 32192 63957 32201
rect 63043 32151 63101 32152
rect 63915 32152 63916 32192
rect 63956 32152 63957 32192
rect 64099 32173 64108 32213
rect 64148 32173 64157 32213
rect 64099 32172 64157 32173
rect 64291 32192 64349 32193
rect 63915 32143 63957 32152
rect 64291 32152 64300 32192
rect 64340 32152 64349 32192
rect 64291 32151 64349 32152
rect 64491 32192 64533 32201
rect 64491 32152 64492 32192
rect 64532 32152 64533 32192
rect 64491 32143 64533 32152
rect 65347 32192 65405 32193
rect 65347 32152 65356 32192
rect 65396 32152 65405 32192
rect 65347 32151 65405 32152
rect 65547 32192 65589 32201
rect 65547 32152 65548 32192
rect 65588 32152 65589 32192
rect 65547 32143 65589 32152
rect 66123 32192 66165 32201
rect 66123 32152 66124 32192
rect 66164 32152 66165 32192
rect 66123 32143 66165 32152
rect 66403 32192 66461 32193
rect 66403 32152 66412 32192
rect 66452 32152 66461 32192
rect 66403 32151 66461 32152
rect 66699 32192 66741 32201
rect 66699 32152 66700 32192
rect 66740 32152 66741 32192
rect 66699 32143 66741 32152
rect 67075 32192 67133 32193
rect 67075 32152 67084 32192
rect 67124 32152 67133 32192
rect 67075 32151 67133 32152
rect 67939 32192 67997 32193
rect 67939 32152 67948 32192
rect 67988 32152 67997 32192
rect 67939 32151 67997 32152
rect 69763 32192 69821 32193
rect 69763 32152 69772 32192
rect 69812 32152 69821 32192
rect 69763 32151 69821 32152
rect 69867 32192 69909 32201
rect 69867 32152 69868 32192
rect 69908 32152 69909 32192
rect 69867 32143 69909 32152
rect 70059 32192 70101 32201
rect 70059 32152 70060 32192
rect 70100 32152 70101 32192
rect 70059 32143 70101 32152
rect 70251 32192 70293 32201
rect 70251 32152 70252 32192
rect 70292 32152 70293 32192
rect 70251 32143 70293 32152
rect 70347 32192 70389 32201
rect 70347 32152 70348 32192
rect 70388 32152 70389 32192
rect 70347 32143 70389 32152
rect 70443 32192 70485 32201
rect 70443 32152 70444 32192
rect 70484 32152 70485 32192
rect 70443 32143 70485 32152
rect 70539 32192 70581 32201
rect 70539 32152 70540 32192
rect 70580 32152 70581 32192
rect 70539 32143 70581 32152
rect 70819 32192 70877 32193
rect 70819 32152 70828 32192
rect 70868 32152 70877 32192
rect 70819 32151 70877 32152
rect 70923 32192 70965 32201
rect 70923 32152 70924 32192
rect 70964 32152 70965 32192
rect 70923 32143 70965 32152
rect 71115 32192 71157 32201
rect 71115 32152 71116 32192
rect 71156 32152 71157 32192
rect 71115 32143 71157 32152
rect 71587 32192 71645 32193
rect 71587 32152 71596 32192
rect 71636 32152 71645 32192
rect 71587 32151 71645 32152
rect 71883 32192 71925 32201
rect 71883 32152 71884 32192
rect 71924 32152 71925 32192
rect 71883 32143 71925 32152
rect 72459 32192 72501 32201
rect 72459 32152 72460 32192
rect 72500 32152 72501 32192
rect 72459 32143 72501 32152
rect 72643 32192 72701 32193
rect 72643 32152 72652 32192
rect 72692 32152 72701 32192
rect 72643 32151 72701 32152
rect 75819 32192 75861 32201
rect 75819 32152 75820 32192
rect 75860 32152 75861 32192
rect 75819 32143 75861 32152
rect 76011 32192 76053 32201
rect 76011 32152 76012 32192
rect 76052 32152 76053 32192
rect 76011 32143 76053 32152
rect 76099 32192 76157 32193
rect 76099 32152 76108 32192
rect 76148 32152 76157 32192
rect 76099 32151 76157 32152
rect 76675 32192 76733 32193
rect 76675 32152 76684 32192
rect 76724 32152 76733 32192
rect 76675 32151 76733 32152
rect 76875 32192 76917 32201
rect 76875 32152 76876 32192
rect 76916 32152 76917 32192
rect 76875 32143 76917 32152
rect 77443 32192 77501 32193
rect 77443 32152 77452 32192
rect 77492 32152 77501 32192
rect 77443 32151 77501 32152
rect 78307 32192 78365 32193
rect 78307 32152 78316 32192
rect 78356 32152 78365 32192
rect 78307 32151 78365 32152
rect 49035 32098 49077 32107
rect 59307 32108 59349 32117
rect 59307 32068 59308 32108
rect 59348 32068 59349 32108
rect 59307 32059 59349 32068
rect 79467 32108 79509 32117
rect 79467 32068 79468 32108
rect 79508 32068 79509 32108
rect 79467 32059 79509 32068
rect 40587 32024 40629 32033
rect 40587 31984 40588 32024
rect 40628 31984 40629 32024
rect 40587 31975 40629 31984
rect 53539 32024 53597 32025
rect 53539 31984 53548 32024
rect 53588 31984 53597 32024
rect 53539 31983 53597 31984
rect 56619 32024 56661 32033
rect 56619 31984 56620 32024
rect 56660 31984 56661 32024
rect 56619 31975 56661 31984
rect 59011 32024 59069 32025
rect 59011 31984 59020 32024
rect 59060 31984 59069 32024
rect 59011 31983 59069 31984
rect 63715 32024 63773 32025
rect 63715 31984 63724 32024
rect 63764 31984 63773 32024
rect 63715 31983 63773 31984
rect 65451 32024 65493 32033
rect 65451 31984 65452 32024
rect 65492 31984 65493 32024
rect 65451 31975 65493 31984
rect 65731 32024 65789 32025
rect 65731 31984 65740 32024
rect 65780 31984 65789 32024
rect 65731 31983 65789 31984
rect 72259 32024 72317 32025
rect 72259 31984 72268 32024
rect 72308 31984 72317 32024
rect 72259 31983 72317 31984
rect 72555 32024 72597 32033
rect 72555 31984 72556 32024
rect 72596 31984 72597 32024
rect 72555 31975 72597 31984
rect 72843 32024 72885 32033
rect 72843 31984 72844 32024
rect 72884 31984 72885 32024
rect 72843 31975 72885 31984
rect 74091 32024 74133 32033
rect 74091 31984 74092 32024
rect 74132 31984 74133 32024
rect 74091 31975 74133 31984
rect 42987 31940 43029 31949
rect 42987 31900 42988 31940
rect 43028 31900 43029 31940
rect 42987 31891 43029 31900
rect 45667 31940 45725 31941
rect 45667 31900 45676 31940
rect 45716 31900 45725 31940
rect 45667 31899 45725 31900
rect 49611 31940 49653 31949
rect 49611 31900 49612 31940
rect 49652 31900 49653 31940
rect 49611 31891 49653 31900
rect 59883 31940 59925 31949
rect 59883 31900 59884 31940
rect 59924 31900 59925 31940
rect 59883 31891 59925 31900
rect 64011 31940 64053 31949
rect 64011 31900 64012 31940
rect 64052 31900 64053 31940
rect 64011 31891 64053 31900
rect 64395 31940 64437 31949
rect 64395 31900 64396 31940
rect 64436 31900 64437 31940
rect 64395 31891 64437 31900
rect 69091 31940 69149 31941
rect 69091 31900 69100 31940
rect 69140 31900 69149 31940
rect 69091 31899 69149 31900
rect 71115 31940 71157 31949
rect 71115 31900 71116 31940
rect 71156 31900 71157 31940
rect 71115 31891 71157 31900
rect 576 31772 79584 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 75112 31772
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75480 31732 79584 31772
rect 576 31708 79584 31732
rect 42691 31604 42749 31605
rect 42691 31564 42700 31604
rect 42740 31564 42749 31604
rect 42691 31563 42749 31564
rect 43947 31604 43989 31613
rect 43947 31564 43948 31604
rect 43988 31564 43989 31604
rect 43947 31555 43989 31564
rect 48843 31604 48885 31613
rect 48843 31564 48844 31604
rect 48884 31564 48885 31604
rect 48843 31555 48885 31564
rect 51147 31604 51189 31613
rect 51147 31564 51148 31604
rect 51188 31564 51189 31604
rect 51147 31555 51189 31564
rect 51819 31604 51861 31613
rect 51819 31564 51820 31604
rect 51860 31564 51861 31604
rect 51819 31555 51861 31564
rect 55171 31604 55229 31605
rect 55171 31564 55180 31604
rect 55220 31564 55229 31604
rect 55171 31563 55229 31564
rect 63051 31604 63093 31613
rect 63051 31564 63052 31604
rect 63092 31564 63093 31604
rect 63051 31555 63093 31564
rect 66411 31604 66453 31613
rect 66411 31564 66412 31604
rect 66452 31564 66453 31604
rect 66411 31555 66453 31564
rect 71115 31604 71157 31613
rect 71115 31564 71116 31604
rect 71156 31564 71157 31604
rect 71115 31555 71157 31564
rect 76003 31604 76061 31605
rect 76003 31564 76012 31604
rect 76052 31564 76061 31604
rect 76003 31563 76061 31564
rect 48363 31520 48405 31529
rect 48363 31480 48364 31520
rect 48404 31480 48405 31520
rect 48363 31471 48405 31480
rect 49707 31520 49749 31529
rect 49707 31480 49708 31520
rect 49748 31480 49749 31520
rect 49707 31471 49749 31480
rect 61131 31520 61173 31529
rect 61131 31480 61132 31520
rect 61172 31480 61173 31520
rect 50947 31478 51005 31479
rect 50947 31438 50956 31478
rect 50996 31438 51005 31478
rect 61131 31471 61173 31480
rect 63627 31520 63669 31529
rect 63627 31480 63628 31520
rect 63668 31480 63669 31520
rect 63627 31471 63669 31480
rect 67275 31520 67317 31529
rect 67275 31480 67276 31520
rect 67316 31480 67317 31520
rect 67275 31471 67317 31480
rect 68811 31520 68853 31529
rect 68811 31480 68812 31520
rect 68852 31480 68853 31520
rect 68811 31471 68853 31480
rect 72267 31520 72309 31529
rect 72267 31480 72268 31520
rect 72308 31480 72309 31520
rect 72267 31471 72309 31480
rect 77835 31520 77877 31529
rect 77835 31480 77836 31520
rect 77876 31480 77877 31520
rect 77835 31471 77877 31480
rect 50947 31437 51005 31438
rect 51619 31436 51677 31437
rect 51619 31396 51628 31436
rect 51668 31396 51677 31436
rect 51619 31395 51677 31396
rect 60643 31436 60701 31437
rect 60643 31396 60652 31436
rect 60692 31396 60701 31436
rect 60643 31395 60701 31396
rect 70915 31436 70973 31437
rect 70915 31396 70924 31436
rect 70964 31396 70973 31436
rect 70915 31395 70973 31396
rect 63357 31363 63399 31372
rect 40483 31352 40541 31353
rect 40483 31312 40492 31352
rect 40532 31312 40541 31352
rect 40483 31311 40541 31312
rect 41347 31352 41405 31353
rect 41347 31312 41356 31352
rect 41396 31312 41405 31352
rect 41347 31311 41405 31312
rect 43083 31352 43125 31361
rect 43083 31312 43084 31352
rect 43124 31312 43125 31352
rect 43083 31303 43125 31312
rect 43363 31352 43421 31353
rect 43363 31312 43372 31352
rect 43412 31312 43421 31352
rect 43363 31311 43421 31312
rect 43651 31352 43709 31353
rect 43651 31312 43660 31352
rect 43700 31312 43709 31352
rect 43651 31311 43709 31312
rect 43755 31352 43797 31361
rect 43755 31312 43756 31352
rect 43796 31312 43797 31352
rect 43755 31303 43797 31312
rect 43947 31352 43989 31361
rect 43947 31312 43948 31352
rect 43988 31312 43989 31352
rect 43947 31303 43989 31312
rect 48547 31352 48605 31353
rect 48547 31312 48556 31352
rect 48596 31312 48605 31352
rect 48547 31311 48605 31312
rect 48651 31352 48693 31361
rect 48651 31312 48652 31352
rect 48692 31312 48693 31352
rect 48651 31303 48693 31312
rect 48843 31352 48885 31361
rect 48843 31312 48844 31352
rect 48884 31312 48885 31352
rect 48843 31303 48885 31312
rect 49227 31352 49269 31361
rect 49227 31312 49228 31352
rect 49268 31312 49269 31352
rect 49227 31303 49269 31312
rect 49419 31352 49461 31361
rect 49419 31312 49420 31352
rect 49460 31312 49461 31352
rect 49419 31303 49461 31312
rect 49507 31352 49565 31353
rect 49507 31312 49516 31352
rect 49556 31312 49565 31352
rect 49507 31311 49565 31312
rect 49707 31352 49749 31361
rect 49707 31312 49708 31352
rect 49748 31312 49749 31352
rect 49707 31303 49749 31312
rect 49899 31352 49941 31361
rect 49899 31312 49900 31352
rect 49940 31312 49941 31352
rect 49899 31303 49941 31312
rect 49987 31352 50045 31353
rect 49987 31312 49996 31352
rect 50036 31312 50045 31352
rect 49987 31311 50045 31312
rect 50275 31352 50333 31353
rect 50275 31312 50284 31352
rect 50324 31312 50333 31352
rect 50275 31311 50333 31312
rect 50571 31352 50613 31361
rect 50571 31312 50572 31352
rect 50612 31312 50613 31352
rect 50571 31303 50613 31312
rect 50667 31352 50709 31361
rect 50667 31312 50668 31352
rect 50708 31312 50709 31352
rect 50667 31303 50709 31312
rect 51147 31352 51189 31361
rect 51147 31312 51148 31352
rect 51188 31312 51189 31352
rect 51147 31303 51189 31312
rect 51339 31352 51381 31361
rect 51339 31312 51340 31352
rect 51380 31312 51381 31352
rect 51339 31303 51381 31312
rect 51427 31352 51485 31353
rect 51427 31312 51436 31352
rect 51476 31312 51485 31352
rect 51427 31311 51485 31312
rect 53155 31352 53213 31353
rect 53155 31312 53164 31352
rect 53204 31312 53213 31352
rect 53155 31311 53213 31312
rect 54019 31352 54077 31353
rect 54019 31312 54028 31352
rect 54068 31312 54077 31352
rect 54019 31311 54077 31312
rect 55555 31352 55613 31353
rect 55555 31312 55564 31352
rect 55604 31312 55613 31352
rect 55555 31311 55613 31312
rect 55755 31352 55797 31361
rect 55755 31312 55756 31352
rect 55796 31312 55797 31352
rect 55755 31303 55797 31312
rect 56515 31352 56573 31353
rect 56515 31312 56524 31352
rect 56564 31312 56573 31352
rect 56515 31311 56573 31312
rect 57379 31352 57437 31353
rect 57379 31312 57388 31352
rect 57428 31312 57437 31352
rect 57379 31311 57437 31312
rect 59595 31352 59637 31361
rect 59595 31312 59596 31352
rect 59636 31312 59637 31352
rect 59595 31303 59637 31312
rect 59787 31352 59829 31361
rect 59787 31312 59788 31352
rect 59828 31312 59829 31352
rect 59787 31303 59829 31312
rect 59875 31352 59933 31353
rect 59875 31312 59884 31352
rect 59924 31312 59933 31352
rect 59875 31311 59933 31312
rect 62571 31352 62613 31361
rect 62571 31312 62572 31352
rect 62612 31312 62613 31352
rect 62571 31303 62613 31312
rect 62763 31352 62805 31361
rect 62763 31312 62764 31352
rect 62804 31312 62805 31352
rect 62763 31303 62805 31312
rect 62851 31352 62909 31353
rect 62851 31312 62860 31352
rect 62900 31312 62909 31352
rect 62851 31311 62909 31312
rect 63051 31352 63093 31361
rect 63051 31312 63052 31352
rect 63092 31312 63093 31352
rect 63051 31303 63093 31312
rect 63243 31352 63285 31361
rect 63243 31312 63244 31352
rect 63284 31312 63285 31352
rect 63357 31323 63358 31363
rect 63398 31323 63399 31363
rect 63357 31314 63399 31323
rect 66411 31352 66453 31361
rect 63243 31303 63285 31312
rect 66411 31312 66412 31352
rect 66452 31312 66453 31352
rect 66411 31303 66453 31312
rect 66603 31352 66645 31361
rect 66603 31312 66604 31352
rect 66644 31312 66645 31352
rect 66603 31303 66645 31312
rect 66691 31352 66749 31353
rect 66691 31312 66700 31352
rect 66740 31312 66749 31352
rect 66691 31311 66749 31312
rect 66883 31352 66941 31353
rect 66883 31312 66892 31352
rect 66932 31312 66941 31352
rect 66883 31311 66941 31312
rect 67083 31352 67125 31361
rect 67083 31312 67084 31352
rect 67124 31312 67125 31352
rect 67083 31303 67125 31312
rect 70539 31352 70581 31361
rect 70539 31312 70540 31352
rect 70580 31312 70581 31352
rect 70539 31303 70581 31312
rect 70635 31352 70677 31361
rect 70635 31312 70636 31352
rect 70676 31312 70677 31352
rect 70635 31303 70677 31312
rect 70731 31352 70773 31361
rect 70731 31312 70732 31352
rect 70772 31312 70773 31352
rect 70731 31303 70773 31312
rect 71395 31352 71453 31353
rect 71395 31312 71404 31352
rect 71444 31312 71453 31352
rect 71395 31311 71453 31312
rect 71595 31352 71637 31361
rect 71595 31312 71596 31352
rect 71636 31312 71637 31352
rect 71595 31303 71637 31312
rect 73987 31352 74045 31353
rect 73987 31312 73996 31352
rect 74036 31312 74045 31352
rect 73987 31311 74045 31312
rect 74851 31352 74909 31353
rect 74851 31312 74860 31352
rect 74900 31312 74909 31352
rect 74851 31311 74909 31312
rect 76971 31352 77013 31361
rect 76971 31312 76972 31352
rect 77012 31312 77013 31352
rect 76971 31303 77013 31312
rect 77155 31352 77213 31353
rect 77155 31312 77164 31352
rect 77204 31312 77213 31352
rect 77155 31311 77213 31312
rect 77443 31352 77501 31353
rect 77443 31312 77452 31352
rect 77492 31312 77501 31352
rect 77443 31311 77501 31312
rect 77643 31352 77685 31361
rect 77643 31312 77644 31352
rect 77684 31312 77685 31352
rect 77643 31303 77685 31312
rect 40107 31268 40149 31277
rect 40107 31228 40108 31268
rect 40148 31228 40149 31268
rect 40107 31219 40149 31228
rect 42987 31268 43029 31277
rect 42987 31228 42988 31268
rect 43028 31228 43029 31268
rect 42987 31219 43029 31228
rect 52779 31268 52821 31277
rect 52779 31228 52780 31268
rect 52820 31228 52821 31268
rect 52779 31219 52821 31228
rect 55659 31268 55701 31277
rect 55659 31228 55660 31268
rect 55700 31228 55701 31268
rect 55659 31219 55701 31228
rect 56139 31268 56181 31277
rect 56139 31228 56140 31268
rect 56180 31228 56181 31268
rect 56139 31219 56181 31228
rect 62667 31268 62709 31277
rect 62667 31228 62668 31268
rect 62708 31228 62709 31268
rect 62667 31219 62709 31228
rect 66987 31268 67029 31277
rect 66987 31228 66988 31268
rect 67028 31228 67029 31268
rect 66987 31219 67029 31228
rect 71499 31268 71541 31277
rect 71499 31228 71500 31268
rect 71540 31228 71541 31268
rect 71499 31219 71541 31228
rect 73611 31268 73653 31277
rect 73611 31228 73612 31268
rect 73652 31228 73653 31268
rect 73611 31219 73653 31228
rect 77067 31268 77109 31277
rect 77067 31228 77068 31268
rect 77108 31228 77109 31268
rect 77067 31219 77109 31228
rect 77547 31268 77589 31277
rect 77547 31228 77548 31268
rect 77588 31228 77589 31268
rect 77547 31219 77589 31228
rect 42499 31184 42557 31185
rect 42499 31144 42508 31184
rect 42548 31144 42557 31184
rect 42499 31143 42557 31144
rect 49315 31184 49373 31185
rect 49315 31144 49324 31184
rect 49364 31144 49373 31184
rect 49315 31143 49373 31144
rect 51819 31184 51861 31193
rect 51819 31144 51820 31184
rect 51860 31144 51861 31184
rect 51819 31135 51861 31144
rect 55171 31184 55229 31185
rect 55171 31144 55180 31184
rect 55220 31144 55229 31184
rect 55171 31143 55229 31144
rect 58531 31184 58589 31185
rect 58531 31144 58540 31184
rect 58580 31144 58589 31184
rect 58531 31143 58589 31144
rect 59683 31184 59741 31185
rect 59683 31144 59692 31184
rect 59732 31144 59741 31184
rect 59683 31143 59741 31144
rect 60459 31184 60501 31193
rect 60459 31144 60460 31184
rect 60500 31144 60501 31184
rect 60459 31135 60501 31144
rect 70435 31184 70493 31185
rect 70435 31144 70444 31184
rect 70484 31144 70493 31184
rect 70435 31143 70493 31144
rect 71115 31184 71157 31193
rect 71115 31144 71116 31184
rect 71156 31144 71157 31184
rect 71115 31135 71157 31144
rect 76003 31184 76061 31185
rect 76003 31144 76012 31184
rect 76052 31144 76061 31184
rect 76003 31143 76061 31144
rect 576 31016 79584 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 76352 31016
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76720 30976 79584 31016
rect 576 30952 79584 30976
rect 40971 30848 41013 30857
rect 40971 30808 40972 30848
rect 41012 30808 41013 30848
rect 40971 30799 41013 30808
rect 52107 30848 52149 30857
rect 52107 30808 52108 30848
rect 52148 30808 52149 30848
rect 52107 30799 52149 30808
rect 56035 30848 56093 30849
rect 56035 30808 56044 30848
rect 56084 30808 56093 30848
rect 56035 30807 56093 30808
rect 60939 30848 60981 30857
rect 60939 30808 60940 30848
rect 60980 30808 60981 30848
rect 60939 30799 60981 30808
rect 61707 30848 61749 30857
rect 61707 30808 61708 30848
rect 61748 30808 61749 30848
rect 61707 30799 61749 30808
rect 62755 30848 62813 30849
rect 62755 30808 62764 30848
rect 62804 30808 62813 30848
rect 62755 30807 62813 30808
rect 75427 30848 75485 30849
rect 75427 30808 75436 30848
rect 75476 30808 75485 30848
rect 75427 30807 75485 30808
rect 43371 30764 43413 30773
rect 43371 30724 43372 30764
rect 43412 30724 43413 30764
rect 43371 30715 43413 30724
rect 48075 30764 48117 30773
rect 48075 30724 48076 30764
rect 48116 30724 48117 30764
rect 48075 30715 48117 30724
rect 50859 30764 50901 30773
rect 50859 30724 50860 30764
rect 50900 30724 50901 30764
rect 50859 30715 50901 30724
rect 55467 30764 55509 30773
rect 55467 30724 55468 30764
rect 55508 30724 55509 30764
rect 55467 30715 55509 30724
rect 57771 30764 57813 30773
rect 57771 30724 57772 30764
rect 57812 30724 57813 30764
rect 57771 30715 57813 30724
rect 71307 30764 71349 30773
rect 71307 30724 71308 30764
rect 71348 30724 71349 30764
rect 71307 30715 71349 30724
rect 74859 30764 74901 30773
rect 74859 30724 74860 30764
rect 74900 30724 74901 30764
rect 74859 30715 74901 30724
rect 66123 30693 66165 30702
rect 59011 30691 59069 30692
rect 42987 30680 43029 30689
rect 42795 30669 42837 30678
rect 42795 30629 42796 30669
rect 42836 30629 42837 30669
rect 42987 30640 42988 30680
rect 43028 30640 43029 30680
rect 42987 30631 43029 30640
rect 43075 30680 43133 30681
rect 43075 30640 43084 30680
rect 43124 30640 43133 30680
rect 43075 30639 43133 30640
rect 43275 30680 43317 30689
rect 43275 30640 43276 30680
rect 43316 30640 43317 30680
rect 43275 30631 43317 30640
rect 43459 30680 43517 30681
rect 43459 30640 43468 30680
rect 43508 30640 43517 30680
rect 43459 30639 43517 30640
rect 43947 30680 43989 30689
rect 43947 30640 43948 30680
rect 43988 30640 43989 30680
rect 43947 30631 43989 30640
rect 44139 30680 44181 30689
rect 44139 30640 44140 30680
rect 44180 30640 44181 30680
rect 44139 30631 44181 30640
rect 44227 30680 44285 30681
rect 44227 30640 44236 30680
rect 44276 30640 44285 30680
rect 44227 30639 44285 30640
rect 44907 30680 44949 30689
rect 44907 30640 44908 30680
rect 44948 30640 44949 30680
rect 44907 30631 44949 30640
rect 45003 30680 45045 30689
rect 45003 30640 45004 30680
rect 45044 30640 45045 30680
rect 45003 30631 45045 30640
rect 45099 30680 45141 30689
rect 45099 30640 45100 30680
rect 45140 30640 45141 30680
rect 45099 30631 45141 30640
rect 45195 30680 45237 30689
rect 45195 30640 45196 30680
rect 45236 30640 45237 30680
rect 45195 30631 45237 30640
rect 45867 30680 45909 30689
rect 45867 30640 45868 30680
rect 45908 30640 45909 30680
rect 45867 30631 45909 30640
rect 46051 30680 46109 30681
rect 46051 30640 46060 30680
rect 46100 30640 46109 30680
rect 46051 30639 46109 30640
rect 46243 30680 46301 30681
rect 46243 30640 46252 30680
rect 46292 30640 46301 30680
rect 46243 30639 46301 30640
rect 46347 30680 46389 30689
rect 46347 30640 46348 30680
rect 46388 30640 46389 30680
rect 46347 30631 46389 30640
rect 46539 30680 46581 30689
rect 46539 30640 46540 30680
rect 46580 30640 46581 30680
rect 46539 30631 46581 30640
rect 48451 30680 48509 30681
rect 48451 30640 48460 30680
rect 48500 30640 48509 30680
rect 48451 30639 48509 30640
rect 49315 30680 49373 30681
rect 49315 30640 49324 30680
rect 49364 30640 49373 30680
rect 49315 30639 49373 30640
rect 50755 30680 50813 30681
rect 50755 30640 50764 30680
rect 50804 30640 50813 30680
rect 50755 30639 50813 30640
rect 50955 30680 50997 30689
rect 50955 30640 50956 30680
rect 50996 30640 50997 30680
rect 50955 30631 50997 30640
rect 51139 30680 51197 30681
rect 51139 30640 51148 30680
rect 51188 30640 51197 30680
rect 51139 30639 51197 30640
rect 51339 30680 51381 30689
rect 51339 30640 51340 30680
rect 51380 30640 51381 30680
rect 51339 30631 51381 30640
rect 54507 30680 54549 30689
rect 54507 30640 54508 30680
rect 54548 30640 54549 30680
rect 54507 30631 54549 30640
rect 54699 30680 54741 30689
rect 54699 30640 54700 30680
rect 54740 30640 54741 30680
rect 54699 30631 54741 30640
rect 54787 30680 54845 30681
rect 54787 30640 54796 30680
rect 54836 30640 54845 30680
rect 54787 30639 54845 30640
rect 55075 30680 55133 30681
rect 55075 30640 55084 30680
rect 55124 30640 55133 30680
rect 55075 30639 55133 30640
rect 55371 30680 55413 30689
rect 55371 30640 55372 30680
rect 55412 30640 55413 30680
rect 55371 30631 55413 30640
rect 55947 30680 55989 30689
rect 55947 30640 55948 30680
rect 55988 30640 55989 30680
rect 55947 30631 55989 30640
rect 56139 30680 56181 30689
rect 56139 30640 56140 30680
rect 56180 30640 56181 30680
rect 56139 30631 56181 30640
rect 56227 30680 56285 30681
rect 56227 30640 56236 30680
rect 56276 30640 56285 30680
rect 56227 30639 56285 30640
rect 56419 30680 56477 30681
rect 56419 30640 56428 30680
rect 56468 30640 56477 30680
rect 56419 30639 56477 30640
rect 56619 30680 56661 30689
rect 56619 30640 56620 30680
rect 56660 30640 56661 30680
rect 56619 30631 56661 30640
rect 58147 30680 58205 30681
rect 58147 30640 58156 30680
rect 58196 30640 58205 30680
rect 59011 30651 59020 30691
rect 59060 30651 59069 30691
rect 59011 30650 59069 30651
rect 61123 30680 61181 30681
rect 58147 30639 58205 30640
rect 61123 30640 61132 30680
rect 61172 30640 61181 30680
rect 61123 30639 61181 30640
rect 61323 30680 61365 30689
rect 61323 30640 61324 30680
rect 61364 30640 61365 30680
rect 61323 30631 61365 30640
rect 62667 30680 62709 30689
rect 62667 30640 62668 30680
rect 62708 30640 62709 30680
rect 62667 30631 62709 30640
rect 62859 30680 62901 30689
rect 62859 30640 62860 30680
rect 62900 30640 62901 30680
rect 62859 30631 62901 30640
rect 62947 30680 63005 30681
rect 62947 30640 62956 30680
rect 62996 30640 63005 30680
rect 62947 30639 63005 30640
rect 63147 30680 63189 30689
rect 63147 30640 63148 30680
rect 63188 30640 63189 30680
rect 63147 30631 63189 30640
rect 63523 30680 63581 30681
rect 63523 30640 63532 30680
rect 63572 30640 63581 30680
rect 63523 30639 63581 30640
rect 64387 30680 64445 30681
rect 64387 30640 64396 30680
rect 64436 30640 64445 30680
rect 64387 30639 64445 30640
rect 65923 30680 65981 30681
rect 65923 30640 65932 30680
rect 65972 30640 65981 30680
rect 66123 30653 66124 30693
rect 66164 30653 66165 30693
rect 66123 30644 66165 30653
rect 68235 30680 68277 30689
rect 65923 30639 65981 30640
rect 68235 30640 68236 30680
rect 68276 30640 68277 30680
rect 68235 30631 68277 30640
rect 68611 30680 68669 30681
rect 68611 30640 68620 30680
rect 68660 30640 68669 30680
rect 68611 30639 68669 30640
rect 69475 30680 69533 30681
rect 69475 30640 69484 30680
rect 69524 30640 69533 30680
rect 69475 30639 69533 30640
rect 70915 30680 70973 30681
rect 70915 30640 70924 30680
rect 70964 30640 70973 30680
rect 70915 30639 70973 30640
rect 71211 30680 71253 30689
rect 71211 30640 71212 30680
rect 71252 30640 71253 30680
rect 71211 30631 71253 30640
rect 71787 30680 71829 30689
rect 71787 30640 71788 30680
rect 71828 30640 71829 30680
rect 71787 30631 71829 30640
rect 72163 30680 72221 30681
rect 72163 30640 72172 30680
rect 72212 30640 72221 30680
rect 72163 30639 72221 30640
rect 73027 30680 73085 30681
rect 73027 30640 73036 30680
rect 73076 30640 73085 30680
rect 73027 30639 73085 30640
rect 74955 30680 74997 30689
rect 74955 30640 74956 30680
rect 74996 30640 74997 30680
rect 74955 30631 74997 30640
rect 75051 30680 75093 30689
rect 75051 30640 75052 30680
rect 75092 30640 75093 30680
rect 75051 30631 75093 30640
rect 75147 30680 75189 30689
rect 75147 30640 75148 30680
rect 75188 30640 75189 30680
rect 75147 30631 75189 30640
rect 75339 30680 75381 30689
rect 75339 30640 75340 30680
rect 75380 30640 75381 30680
rect 75339 30631 75381 30640
rect 75531 30680 75573 30689
rect 75531 30640 75532 30680
rect 75572 30640 75573 30680
rect 75531 30631 75573 30640
rect 75619 30680 75677 30681
rect 75619 30640 75628 30680
rect 75668 30640 75677 30680
rect 75619 30639 75677 30640
rect 76195 30680 76253 30681
rect 76195 30640 76204 30680
rect 76244 30640 76253 30680
rect 76195 30639 76253 30640
rect 76491 30680 76533 30689
rect 76491 30640 76492 30680
rect 76532 30640 76533 30680
rect 76491 30631 76533 30640
rect 76587 30680 76629 30689
rect 76587 30640 76588 30680
rect 76628 30640 76629 30680
rect 76587 30631 76629 30640
rect 77067 30680 77109 30689
rect 77067 30640 77068 30680
rect 77108 30640 77109 30680
rect 77067 30631 77109 30640
rect 77443 30680 77501 30681
rect 77443 30640 77452 30680
rect 77492 30640 77501 30680
rect 77443 30639 77501 30640
rect 78307 30680 78365 30681
rect 78307 30640 78316 30680
rect 78356 30640 78365 30680
rect 78307 30639 78365 30640
rect 42795 30620 42837 30629
rect 40579 30596 40637 30597
rect 40579 30556 40588 30596
rect 40628 30556 40637 30596
rect 40579 30555 40637 30556
rect 41155 30596 41213 30597
rect 41155 30556 41164 30596
rect 41204 30556 41213 30596
rect 41155 30555 41213 30556
rect 42403 30596 42461 30597
rect 42403 30556 42412 30596
rect 42452 30556 42461 30596
rect 42403 30555 42461 30556
rect 51523 30596 51581 30597
rect 51523 30556 51532 30596
rect 51572 30556 51581 30596
rect 51523 30555 51581 30556
rect 51907 30596 51965 30597
rect 51907 30556 51916 30596
rect 51956 30556 51965 30596
rect 56523 30596 56565 30605
rect 51907 30555 51965 30556
rect 53259 30554 53301 30563
rect 43947 30512 43989 30521
rect 43947 30472 43948 30512
rect 43988 30472 43989 30512
rect 43947 30463 43989 30472
rect 44427 30512 44469 30521
rect 44427 30472 44428 30512
rect 44468 30472 44469 30512
rect 44427 30463 44469 30472
rect 47019 30512 47061 30521
rect 47019 30472 47020 30512
rect 47060 30472 47061 30512
rect 47019 30463 47061 30472
rect 52299 30512 52341 30521
rect 52299 30472 52300 30512
rect 52340 30472 52341 30512
rect 53259 30514 53260 30554
rect 53300 30514 53301 30554
rect 56523 30556 56524 30596
rect 56564 30556 56565 30596
rect 56523 30547 56565 30556
rect 60547 30596 60605 30597
rect 60547 30556 60556 30596
rect 60596 30556 60605 30596
rect 60547 30555 60605 30556
rect 60739 30596 60797 30597
rect 60739 30556 60748 30596
rect 60788 30556 60797 30596
rect 60739 30555 60797 30556
rect 61507 30596 61565 30597
rect 61507 30556 61516 30596
rect 61556 30556 61565 30596
rect 61507 30555 61565 30556
rect 53259 30505 53301 30514
rect 54507 30512 54549 30521
rect 52299 30463 52341 30472
rect 54507 30472 54508 30512
rect 54548 30472 54549 30512
rect 54507 30463 54549 30472
rect 55747 30512 55805 30513
rect 55747 30472 55756 30512
rect 55796 30472 55805 30512
rect 55747 30471 55805 30472
rect 66507 30512 66549 30521
rect 66507 30472 66508 30512
rect 66548 30472 66549 30512
rect 66507 30463 66549 30472
rect 71587 30512 71645 30513
rect 71587 30472 71596 30512
rect 71636 30472 71645 30512
rect 71587 30471 71645 30472
rect 76867 30512 76925 30513
rect 76867 30472 76876 30512
rect 76916 30472 76925 30512
rect 76867 30471 76925 30472
rect 79459 30512 79517 30513
rect 79459 30472 79468 30512
rect 79508 30472 79517 30512
rect 79459 30471 79517 30472
rect 40779 30428 40821 30437
rect 40779 30388 40780 30428
rect 40820 30388 40821 30428
rect 40779 30379 40821 30388
rect 40971 30428 41013 30437
rect 40971 30388 40972 30428
rect 41012 30388 41013 30428
rect 40971 30379 41013 30388
rect 42603 30428 42645 30437
rect 42603 30388 42604 30428
rect 42644 30388 42645 30428
rect 42603 30379 42645 30388
rect 42795 30428 42837 30437
rect 42795 30388 42796 30428
rect 42836 30388 42837 30428
rect 42795 30379 42837 30388
rect 45963 30428 46005 30437
rect 45963 30388 45964 30428
rect 46004 30388 46005 30428
rect 45963 30379 46005 30388
rect 46539 30428 46581 30437
rect 46539 30388 46540 30428
rect 46580 30388 46581 30428
rect 46539 30379 46581 30388
rect 50467 30428 50525 30429
rect 50467 30388 50476 30428
rect 50516 30388 50525 30428
rect 50467 30387 50525 30388
rect 51243 30428 51285 30437
rect 51243 30388 51244 30428
rect 51284 30388 51285 30428
rect 51243 30379 51285 30388
rect 51723 30428 51765 30437
rect 51723 30388 51724 30428
rect 51764 30388 51765 30428
rect 51723 30379 51765 30388
rect 52107 30428 52149 30437
rect 52107 30388 52108 30428
rect 52148 30388 52149 30428
rect 52107 30379 52149 30388
rect 60163 30428 60221 30429
rect 60163 30388 60172 30428
rect 60212 30388 60221 30428
rect 60163 30387 60221 30388
rect 60363 30428 60405 30437
rect 60363 30388 60364 30428
rect 60404 30388 60405 30428
rect 60363 30379 60405 30388
rect 60939 30428 60981 30437
rect 60939 30388 60940 30428
rect 60980 30388 60981 30428
rect 60939 30379 60981 30388
rect 61227 30428 61269 30437
rect 61227 30388 61228 30428
rect 61268 30388 61269 30428
rect 61227 30379 61269 30388
rect 61707 30428 61749 30437
rect 61707 30388 61708 30428
rect 61748 30388 61749 30428
rect 61707 30379 61749 30388
rect 65539 30428 65597 30429
rect 65539 30388 65548 30428
rect 65588 30388 65597 30428
rect 65539 30387 65597 30388
rect 66027 30428 66069 30437
rect 66027 30388 66028 30428
rect 66068 30388 66069 30428
rect 66027 30379 66069 30388
rect 70627 30428 70685 30429
rect 70627 30388 70636 30428
rect 70676 30388 70685 30428
rect 70627 30387 70685 30388
rect 74179 30428 74237 30429
rect 74179 30388 74188 30428
rect 74228 30388 74237 30428
rect 74179 30387 74237 30388
rect 576 30260 79584 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 75112 30260
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75480 30220 79584 30260
rect 576 30196 79584 30220
rect 40587 30092 40629 30101
rect 40587 30052 40588 30092
rect 40628 30052 40629 30092
rect 40587 30043 40629 30052
rect 45955 30092 46013 30093
rect 45955 30052 45964 30092
rect 46004 30052 46013 30092
rect 45955 30051 46013 30052
rect 46251 30092 46293 30101
rect 46251 30052 46252 30092
rect 46292 30052 46293 30092
rect 46251 30043 46293 30052
rect 50947 30092 51005 30093
rect 50947 30052 50956 30092
rect 50996 30052 51005 30092
rect 50947 30051 51005 30052
rect 54795 30092 54837 30101
rect 54795 30052 54796 30092
rect 54836 30052 54837 30092
rect 54795 30043 54837 30052
rect 56427 30092 56469 30101
rect 56427 30052 56428 30092
rect 56468 30052 56469 30092
rect 56427 30043 56469 30052
rect 58827 30092 58869 30101
rect 58827 30052 58828 30092
rect 58868 30052 58869 30092
rect 58827 30043 58869 30052
rect 63723 30092 63765 30101
rect 63723 30052 63724 30092
rect 63764 30052 63765 30092
rect 63723 30043 63765 30052
rect 69099 30092 69141 30101
rect 69099 30052 69100 30092
rect 69140 30052 69141 30092
rect 69099 30043 69141 30052
rect 69675 30092 69717 30101
rect 69675 30052 69676 30092
rect 69716 30052 69717 30092
rect 69675 30043 69717 30052
rect 71499 30092 71541 30101
rect 71499 30052 71500 30092
rect 71540 30052 71541 30092
rect 71499 30043 71541 30052
rect 75723 30092 75765 30101
rect 75723 30052 75724 30092
rect 75764 30052 75765 30092
rect 75723 30043 75765 30052
rect 77067 30092 77109 30101
rect 77067 30052 77068 30092
rect 77108 30052 77109 30092
rect 77067 30043 77109 30052
rect 38955 30008 38997 30017
rect 38955 29968 38956 30008
rect 38996 29968 38997 30008
rect 38955 29959 38997 29968
rect 42315 30008 42357 30017
rect 42315 29968 42316 30008
rect 42356 29968 42357 30008
rect 42315 29959 42357 29968
rect 55755 30008 55797 30017
rect 55755 29968 55756 30008
rect 55796 29968 55797 30008
rect 55755 29959 55797 29968
rect 56619 30008 56661 30017
rect 56619 29968 56620 30008
rect 56660 29968 56661 30008
rect 56619 29959 56661 29968
rect 58251 30008 58293 30017
rect 58251 29968 58252 30008
rect 58292 29968 58293 30008
rect 58251 29959 58293 29968
rect 60451 30008 60509 30009
rect 60451 29968 60460 30008
rect 60500 29968 60509 30008
rect 60451 29967 60509 29968
rect 65059 30008 65117 30009
rect 65059 29968 65068 30008
rect 65108 29968 65117 30008
rect 65059 29967 65117 29968
rect 70347 30008 70389 30017
rect 70347 29968 70348 30008
rect 70388 29968 70389 30008
rect 70347 29959 70389 29968
rect 73899 30008 73941 30017
rect 73899 29968 73900 30008
rect 73940 29968 73941 30008
rect 73899 29959 73941 29968
rect 76587 30008 76629 30017
rect 76587 29968 76588 30008
rect 76628 29968 76629 30008
rect 76587 29959 76629 29968
rect 77547 30008 77589 30017
rect 77547 29968 77548 30008
rect 77588 29968 77589 30008
rect 77547 29959 77589 29968
rect 40003 29924 40061 29925
rect 40003 29884 40012 29924
rect 40052 29884 40061 29924
rect 40003 29883 40061 29884
rect 40387 29924 40445 29925
rect 40387 29884 40396 29924
rect 40436 29884 40445 29924
rect 40387 29883 40445 29884
rect 42115 29924 42173 29925
rect 42115 29884 42124 29924
rect 42164 29884 42173 29924
rect 42115 29883 42173 29884
rect 49315 29924 49373 29925
rect 49315 29884 49324 29924
rect 49364 29884 49373 29924
rect 49315 29883 49373 29884
rect 56227 29924 56285 29925
rect 56227 29884 56236 29924
rect 56276 29884 56285 29924
rect 69283 29924 69341 29925
rect 56227 29883 56285 29884
rect 59011 29911 59069 29912
rect 59011 29871 59020 29911
rect 59060 29871 59069 29911
rect 69283 29884 69292 29924
rect 69332 29884 69341 29924
rect 69283 29883 69341 29884
rect 69475 29924 69533 29925
rect 69475 29884 69484 29924
rect 69524 29884 69533 29924
rect 69475 29883 69533 29884
rect 75043 29924 75101 29925
rect 75043 29884 75052 29924
rect 75092 29884 75101 29924
rect 75043 29883 75101 29884
rect 59011 29870 59069 29871
rect 63331 29882 63389 29883
rect 40779 29840 40821 29849
rect 40779 29800 40780 29840
rect 40820 29800 40821 29840
rect 40779 29791 40821 29800
rect 40875 29840 40917 29849
rect 40875 29800 40876 29840
rect 40916 29800 40917 29840
rect 40875 29791 40917 29800
rect 40971 29840 41013 29849
rect 40971 29800 40972 29840
rect 41012 29800 41013 29840
rect 40971 29791 41013 29800
rect 41259 29840 41301 29849
rect 41259 29800 41260 29840
rect 41300 29800 41301 29840
rect 41259 29791 41301 29800
rect 41443 29840 41501 29841
rect 41443 29800 41452 29840
rect 41492 29800 41501 29840
rect 41443 29799 41501 29800
rect 41643 29840 41685 29849
rect 41643 29800 41644 29840
rect 41684 29800 41685 29840
rect 41643 29791 41685 29800
rect 41835 29840 41877 29849
rect 41835 29800 41836 29840
rect 41876 29800 41877 29840
rect 41835 29791 41877 29800
rect 41923 29840 41981 29841
rect 41923 29800 41932 29840
rect 41972 29800 41981 29840
rect 41923 29799 41981 29800
rect 43939 29840 43997 29841
rect 43939 29800 43948 29840
rect 43988 29800 43997 29840
rect 43939 29799 43997 29800
rect 44803 29840 44861 29841
rect 44803 29800 44812 29840
rect 44852 29800 44861 29840
rect 44803 29799 44861 29800
rect 46147 29840 46205 29841
rect 46147 29800 46156 29840
rect 46196 29800 46205 29840
rect 46147 29799 46205 29800
rect 46347 29840 46389 29849
rect 46347 29800 46348 29840
rect 46388 29800 46389 29840
rect 46347 29791 46389 29800
rect 46539 29840 46581 29849
rect 46539 29800 46540 29840
rect 46580 29800 46581 29840
rect 46539 29791 46581 29800
rect 46915 29840 46973 29841
rect 46915 29800 46924 29840
rect 46964 29800 46973 29840
rect 46915 29799 46973 29800
rect 47779 29840 47837 29841
rect 47779 29800 47788 29840
rect 47828 29800 47837 29840
rect 47779 29799 47837 29800
rect 49707 29840 49749 29849
rect 49707 29800 49708 29840
rect 49748 29800 49749 29840
rect 49707 29791 49749 29800
rect 49803 29840 49845 29849
rect 49803 29800 49804 29840
rect 49844 29800 49845 29840
rect 49995 29840 50037 29849
rect 49803 29791 49845 29800
rect 49899 29819 49941 29828
rect 49899 29779 49900 29819
rect 49940 29779 49941 29819
rect 49995 29800 49996 29840
rect 50036 29800 50037 29840
rect 49995 29791 50037 29800
rect 50275 29840 50333 29841
rect 50275 29800 50284 29840
rect 50324 29800 50333 29840
rect 50275 29799 50333 29800
rect 50571 29840 50613 29849
rect 50571 29800 50572 29840
rect 50612 29800 50613 29840
rect 50571 29791 50613 29800
rect 50667 29840 50709 29849
rect 50667 29800 50668 29840
rect 50708 29800 50709 29840
rect 50667 29791 50709 29800
rect 51619 29840 51677 29841
rect 51619 29800 51628 29840
rect 51668 29800 51677 29840
rect 51619 29799 51677 29800
rect 52483 29840 52541 29841
rect 52483 29800 52492 29840
rect 52532 29800 52541 29840
rect 52483 29799 52541 29800
rect 54795 29840 54837 29849
rect 54795 29800 54796 29840
rect 54836 29800 54837 29840
rect 54795 29791 54837 29800
rect 54987 29840 55029 29849
rect 54987 29800 54988 29840
rect 55028 29800 55029 29840
rect 54987 29791 55029 29800
rect 55075 29840 55133 29841
rect 55075 29800 55084 29840
rect 55124 29800 55133 29840
rect 55075 29799 55133 29800
rect 55651 29840 55709 29841
rect 55651 29800 55660 29840
rect 55700 29800 55709 29840
rect 55651 29799 55709 29800
rect 55851 29840 55893 29849
rect 55851 29800 55852 29840
rect 55892 29800 55893 29840
rect 55851 29791 55893 29800
rect 59211 29840 59253 29849
rect 59211 29800 59212 29840
rect 59252 29800 59253 29840
rect 59211 29791 59253 29800
rect 59307 29840 59349 29849
rect 59307 29800 59308 29840
rect 59348 29800 59349 29840
rect 59307 29791 59349 29800
rect 59403 29840 59445 29849
rect 59403 29800 59404 29840
rect 59444 29800 59445 29840
rect 59403 29791 59445 29800
rect 59499 29840 59541 29849
rect 59499 29800 59500 29840
rect 59540 29800 59541 29840
rect 59499 29791 59541 29800
rect 59779 29840 59837 29841
rect 59779 29800 59788 29840
rect 59828 29800 59837 29840
rect 59779 29799 59837 29800
rect 60075 29840 60117 29849
rect 60075 29800 60076 29840
rect 60116 29800 60117 29840
rect 60075 29791 60117 29800
rect 60171 29840 60213 29849
rect 60171 29800 60172 29840
rect 60212 29800 60213 29840
rect 60171 29791 60213 29800
rect 61027 29840 61085 29841
rect 61027 29800 61036 29840
rect 61076 29800 61085 29840
rect 61027 29799 61085 29800
rect 61891 29840 61949 29841
rect 61891 29800 61900 29840
rect 61940 29800 61949 29840
rect 61891 29799 61949 29800
rect 63243 29840 63285 29849
rect 63331 29842 63340 29882
rect 63380 29842 63389 29882
rect 63331 29841 63389 29842
rect 63243 29800 63244 29840
rect 63284 29800 63285 29840
rect 63243 29791 63285 29800
rect 63435 29840 63477 29849
rect 63435 29800 63436 29840
rect 63476 29800 63477 29840
rect 63435 29791 63477 29800
rect 63531 29840 63573 29849
rect 63531 29800 63532 29840
rect 63572 29800 63573 29840
rect 63531 29791 63573 29800
rect 63723 29840 63765 29849
rect 63723 29800 63724 29840
rect 63764 29800 63765 29840
rect 63723 29791 63765 29800
rect 63915 29840 63957 29849
rect 63915 29800 63916 29840
rect 63956 29800 63957 29840
rect 63915 29791 63957 29800
rect 64003 29840 64061 29841
rect 64003 29800 64012 29840
rect 64052 29800 64061 29840
rect 64003 29799 64061 29800
rect 64675 29840 64733 29841
rect 64675 29800 64684 29840
rect 64724 29800 64733 29840
rect 64675 29799 64733 29800
rect 64875 29840 64917 29849
rect 64875 29800 64876 29840
rect 64916 29800 64917 29840
rect 64875 29791 64917 29800
rect 65355 29840 65397 29849
rect 65355 29800 65356 29840
rect 65396 29800 65397 29840
rect 65355 29791 65397 29800
rect 65451 29840 65493 29849
rect 65451 29800 65452 29840
rect 65492 29800 65493 29840
rect 65451 29791 65493 29800
rect 65731 29840 65789 29841
rect 65731 29800 65740 29840
rect 65780 29800 65789 29840
rect 65731 29799 65789 29800
rect 66403 29840 66461 29841
rect 66403 29800 66412 29840
rect 66452 29800 66461 29840
rect 66403 29799 66461 29800
rect 67267 29840 67325 29841
rect 67267 29800 67276 29840
rect 67316 29800 67325 29840
rect 67267 29799 67325 29800
rect 69867 29840 69909 29849
rect 69867 29800 69868 29840
rect 69908 29800 69909 29840
rect 69867 29791 69909 29800
rect 70059 29840 70101 29849
rect 70059 29800 70060 29840
rect 70100 29800 70101 29840
rect 70059 29791 70101 29800
rect 70147 29840 70205 29841
rect 70147 29800 70156 29840
rect 70196 29800 70205 29840
rect 70147 29799 70205 29800
rect 70347 29840 70389 29849
rect 70347 29800 70348 29840
rect 70388 29800 70389 29840
rect 70347 29791 70389 29800
rect 70539 29840 70581 29849
rect 70539 29800 70540 29840
rect 70580 29800 70581 29840
rect 70539 29791 70581 29800
rect 70627 29840 70685 29841
rect 70627 29800 70636 29840
rect 70676 29800 70685 29840
rect 70627 29799 70685 29800
rect 70827 29840 70869 29849
rect 70827 29800 70828 29840
rect 70868 29800 70869 29840
rect 70827 29791 70869 29800
rect 71019 29840 71061 29849
rect 71019 29800 71020 29840
rect 71060 29800 71061 29840
rect 71019 29791 71061 29800
rect 71107 29840 71165 29841
rect 71107 29800 71116 29840
rect 71156 29800 71165 29840
rect 71107 29799 71165 29800
rect 71499 29840 71541 29849
rect 71499 29800 71500 29840
rect 71540 29800 71541 29840
rect 71499 29791 71541 29800
rect 71691 29840 71733 29849
rect 71691 29800 71692 29840
rect 71732 29800 71733 29840
rect 71691 29791 71733 29800
rect 71779 29840 71837 29841
rect 71779 29800 71788 29840
rect 71828 29800 71837 29840
rect 71779 29799 71837 29800
rect 71971 29840 72029 29841
rect 71971 29800 71980 29840
rect 72020 29800 72029 29840
rect 71971 29799 72029 29800
rect 72075 29840 72117 29849
rect 72075 29800 72076 29840
rect 72116 29800 72117 29840
rect 72075 29791 72117 29800
rect 72171 29840 72213 29849
rect 72171 29800 72172 29840
rect 72212 29800 72213 29840
rect 72171 29791 72213 29800
rect 75339 29840 75381 29849
rect 75339 29800 75340 29840
rect 75380 29800 75381 29840
rect 75339 29791 75381 29800
rect 75435 29840 75477 29849
rect 75435 29800 75436 29840
rect 75476 29800 75477 29840
rect 75435 29791 75477 29800
rect 75531 29840 75573 29849
rect 75531 29800 75532 29840
rect 75572 29800 75573 29840
rect 75531 29791 75573 29800
rect 75723 29840 75765 29849
rect 75723 29800 75724 29840
rect 75764 29800 75765 29840
rect 76003 29840 76061 29841
rect 75723 29791 75765 29800
rect 75915 29798 75957 29807
rect 76003 29800 76012 29840
rect 76052 29800 76061 29840
rect 76003 29799 76061 29800
rect 76483 29840 76541 29841
rect 76483 29800 76492 29840
rect 76532 29800 76541 29840
rect 76483 29799 76541 29800
rect 76683 29840 76725 29849
rect 76683 29800 76684 29840
rect 76724 29800 76725 29840
rect 49899 29770 49941 29779
rect 41355 29756 41397 29765
rect 41355 29716 41356 29756
rect 41396 29716 41397 29756
rect 41355 29707 41397 29716
rect 43563 29756 43605 29765
rect 43563 29716 43564 29756
rect 43604 29716 43605 29756
rect 43563 29707 43605 29716
rect 51243 29756 51285 29765
rect 51243 29716 51244 29756
rect 51284 29716 51285 29756
rect 51243 29707 51285 29716
rect 60651 29756 60693 29765
rect 60651 29716 60652 29756
rect 60692 29716 60693 29756
rect 60651 29707 60693 29716
rect 64779 29756 64821 29765
rect 64779 29716 64780 29756
rect 64820 29716 64821 29756
rect 64779 29707 64821 29716
rect 66027 29756 66069 29765
rect 66027 29716 66028 29756
rect 66068 29716 66069 29756
rect 66027 29707 66069 29716
rect 70923 29756 70965 29765
rect 70923 29716 70924 29756
rect 70964 29716 70965 29756
rect 75915 29758 75916 29798
rect 75956 29758 75957 29798
rect 76683 29791 76725 29800
rect 77067 29840 77109 29849
rect 77067 29800 77068 29840
rect 77108 29800 77109 29840
rect 77067 29791 77109 29800
rect 77259 29840 77301 29849
rect 77259 29800 77260 29840
rect 77300 29800 77301 29840
rect 77259 29791 77301 29800
rect 77347 29840 77405 29841
rect 77347 29800 77356 29840
rect 77396 29800 77405 29840
rect 77347 29799 77405 29800
rect 75915 29749 75957 29758
rect 70923 29707 70965 29716
rect 40203 29672 40245 29681
rect 40203 29632 40204 29672
rect 40244 29632 40245 29672
rect 40203 29623 40245 29632
rect 41059 29672 41117 29673
rect 41059 29632 41068 29672
rect 41108 29632 41117 29672
rect 41059 29631 41117 29632
rect 41731 29672 41789 29673
rect 41731 29632 41740 29672
rect 41780 29632 41789 29672
rect 41731 29631 41789 29632
rect 45955 29672 46013 29673
rect 45955 29632 45964 29672
rect 46004 29632 46013 29672
rect 45955 29631 46013 29632
rect 48931 29672 48989 29673
rect 48931 29632 48940 29672
rect 48980 29632 48989 29672
rect 48931 29631 48989 29632
rect 49515 29672 49557 29681
rect 49515 29632 49516 29672
rect 49556 29632 49557 29672
rect 49515 29623 49557 29632
rect 53635 29672 53693 29673
rect 53635 29632 53644 29672
rect 53684 29632 53693 29672
rect 53635 29631 53693 29632
rect 63043 29672 63101 29673
rect 63043 29632 63052 29672
rect 63092 29632 63101 29672
rect 63043 29631 63101 29632
rect 68419 29672 68477 29673
rect 68419 29632 68428 29672
rect 68468 29632 68477 29672
rect 68419 29631 68477 29632
rect 69675 29672 69717 29681
rect 69675 29632 69676 29672
rect 69716 29632 69717 29672
rect 69675 29623 69717 29632
rect 69955 29672 70013 29673
rect 69955 29632 69964 29672
rect 70004 29632 70013 29672
rect 69955 29631 70013 29632
rect 74859 29672 74901 29681
rect 74859 29632 74860 29672
rect 74900 29632 74901 29672
rect 74859 29623 74901 29632
rect 75235 29672 75293 29673
rect 75235 29632 75244 29672
rect 75284 29632 75293 29672
rect 75235 29631 75293 29632
rect 576 29504 79584 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 76352 29504
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76720 29464 79584 29504
rect 576 29440 79584 29464
rect 49611 29336 49653 29345
rect 49611 29296 49612 29336
rect 49652 29296 49653 29336
rect 49611 29287 49653 29296
rect 51043 29336 51101 29337
rect 51043 29296 51052 29336
rect 51092 29296 51101 29336
rect 51043 29295 51101 29296
rect 55267 29336 55325 29337
rect 55267 29296 55276 29336
rect 55316 29296 55325 29336
rect 55267 29295 55325 29296
rect 60451 29336 60509 29337
rect 60451 29296 60460 29336
rect 60500 29296 60509 29336
rect 60451 29295 60509 29296
rect 63427 29336 63485 29337
rect 63427 29296 63436 29336
rect 63476 29296 63485 29336
rect 63427 29295 63485 29296
rect 70243 29336 70301 29337
rect 70243 29296 70252 29336
rect 70292 29296 70301 29336
rect 70243 29295 70301 29296
rect 70731 29336 70773 29345
rect 70731 29296 70732 29336
rect 70772 29296 70773 29336
rect 70731 29287 70773 29296
rect 71691 29336 71733 29345
rect 71691 29296 71692 29336
rect 71732 29296 71733 29336
rect 71691 29287 71733 29296
rect 75811 29336 75869 29337
rect 75811 29296 75820 29336
rect 75860 29296 75869 29336
rect 75811 29295 75869 29296
rect 45963 29252 46005 29261
rect 45963 29212 45964 29252
rect 46004 29212 46005 29252
rect 45963 29203 46005 29212
rect 60939 29252 60981 29261
rect 60939 29212 60940 29252
rect 60980 29212 60981 29252
rect 60939 29203 60981 29212
rect 65739 29252 65781 29261
rect 65739 29212 65740 29252
rect 65780 29212 65781 29252
rect 65739 29203 65781 29212
rect 67659 29252 67701 29261
rect 67659 29212 67660 29252
rect 67700 29212 67701 29252
rect 67659 29203 67701 29212
rect 76491 29252 76533 29261
rect 76491 29212 76492 29252
rect 76532 29212 76533 29252
rect 76491 29203 76533 29212
rect 38475 29168 38517 29177
rect 38475 29128 38476 29168
rect 38516 29128 38517 29168
rect 38475 29119 38517 29128
rect 38851 29168 38909 29169
rect 38851 29128 38860 29168
rect 38900 29128 38909 29168
rect 38851 29127 38909 29128
rect 39715 29168 39773 29169
rect 39715 29128 39724 29168
rect 39764 29128 39773 29168
rect 39715 29127 39773 29128
rect 41355 29168 41397 29177
rect 41355 29128 41356 29168
rect 41396 29128 41397 29168
rect 41355 29119 41397 29128
rect 41451 29168 41493 29177
rect 41451 29128 41452 29168
rect 41492 29128 41493 29168
rect 41451 29119 41493 29128
rect 41731 29168 41789 29169
rect 41731 29128 41740 29168
rect 41780 29128 41789 29168
rect 41731 29127 41789 29128
rect 42019 29168 42077 29169
rect 42019 29128 42028 29168
rect 42068 29128 42077 29168
rect 42019 29127 42077 29128
rect 42123 29168 42165 29177
rect 42123 29128 42124 29168
rect 42164 29128 42165 29168
rect 42123 29119 42165 29128
rect 42315 29168 42357 29177
rect 42315 29128 42316 29168
rect 42356 29128 42357 29168
rect 42315 29119 42357 29128
rect 45099 29168 45141 29177
rect 45099 29128 45100 29168
rect 45140 29128 45141 29168
rect 45099 29119 45141 29128
rect 45291 29168 45333 29177
rect 45291 29128 45292 29168
rect 45332 29128 45333 29168
rect 45291 29119 45333 29128
rect 45379 29168 45437 29169
rect 45379 29128 45388 29168
rect 45428 29128 45437 29168
rect 45379 29127 45437 29128
rect 46059 29168 46101 29177
rect 46059 29128 46060 29168
rect 46100 29128 46101 29168
rect 46059 29119 46101 29128
rect 46339 29168 46397 29169
rect 46339 29128 46348 29168
rect 46388 29128 46397 29168
rect 46339 29127 46397 29128
rect 50187 29168 50229 29177
rect 50187 29128 50188 29168
rect 50228 29128 50229 29168
rect 50187 29119 50229 29128
rect 50379 29168 50421 29177
rect 50379 29128 50380 29168
rect 50420 29128 50421 29168
rect 50379 29119 50421 29128
rect 50467 29168 50525 29169
rect 50467 29128 50476 29168
rect 50516 29128 50525 29168
rect 50467 29127 50525 29128
rect 50851 29168 50909 29169
rect 50851 29128 50860 29168
rect 50900 29128 50909 29168
rect 50851 29127 50909 29128
rect 50955 29168 50997 29177
rect 50955 29128 50956 29168
rect 50996 29128 50997 29168
rect 50955 29119 50997 29128
rect 51147 29168 51189 29177
rect 51147 29128 51148 29168
rect 51188 29128 51189 29168
rect 51147 29119 51189 29128
rect 52875 29168 52917 29177
rect 52875 29128 52876 29168
rect 52916 29128 52917 29168
rect 54115 29168 54173 29169
rect 52875 29119 52917 29128
rect 53251 29132 53309 29133
rect 53251 29092 53260 29132
rect 53300 29092 53309 29132
rect 54115 29128 54124 29168
rect 54164 29128 54173 29168
rect 54115 29127 54173 29128
rect 55467 29168 55509 29177
rect 55467 29128 55468 29168
rect 55508 29128 55509 29168
rect 55467 29119 55509 29128
rect 55563 29168 55605 29177
rect 55563 29128 55564 29168
rect 55604 29128 55605 29168
rect 55563 29119 55605 29128
rect 55659 29168 55701 29177
rect 55659 29128 55660 29168
rect 55700 29128 55701 29168
rect 55659 29119 55701 29128
rect 55755 29168 55797 29177
rect 55755 29128 55756 29168
rect 55796 29128 55797 29168
rect 55755 29119 55797 29128
rect 56139 29168 56181 29177
rect 56139 29128 56140 29168
rect 56180 29128 56181 29168
rect 56139 29119 56181 29128
rect 56515 29168 56573 29169
rect 56515 29128 56524 29168
rect 56564 29128 56573 29168
rect 56515 29127 56573 29128
rect 57379 29168 57437 29169
rect 57379 29128 57388 29168
rect 57428 29128 57437 29168
rect 57379 29127 57437 29128
rect 59587 29168 59645 29169
rect 59587 29128 59596 29168
rect 59636 29128 59645 29168
rect 59587 29127 59645 29128
rect 59691 29168 59733 29177
rect 59691 29128 59692 29168
rect 59732 29128 59733 29168
rect 59691 29119 59733 29128
rect 59883 29168 59925 29177
rect 59883 29128 59884 29168
rect 59924 29128 59925 29168
rect 59883 29119 59925 29128
rect 60363 29168 60405 29177
rect 60363 29128 60364 29168
rect 60404 29128 60405 29168
rect 60363 29119 60405 29128
rect 60555 29168 60597 29177
rect 60555 29128 60556 29168
rect 60596 29128 60597 29168
rect 60555 29119 60597 29128
rect 60643 29168 60701 29169
rect 60643 29128 60652 29168
rect 60692 29128 60701 29168
rect 60643 29127 60701 29128
rect 60843 29168 60885 29177
rect 60843 29128 60844 29168
rect 60884 29128 60885 29168
rect 60843 29119 60885 29128
rect 61027 29168 61085 29169
rect 61027 29128 61036 29168
rect 61076 29128 61085 29168
rect 63531 29168 63573 29177
rect 61027 29127 61085 29128
rect 63339 29157 63381 29166
rect 63339 29117 63340 29157
rect 63380 29117 63381 29157
rect 63531 29128 63532 29168
rect 63572 29128 63573 29168
rect 63531 29119 63573 29128
rect 63619 29168 63677 29169
rect 63619 29128 63628 29168
rect 63668 29128 63677 29168
rect 63619 29127 63677 29128
rect 63819 29168 63861 29177
rect 63819 29128 63820 29168
rect 63860 29128 63861 29168
rect 63819 29119 63861 29128
rect 63915 29168 63957 29177
rect 63915 29128 63916 29168
rect 63956 29128 63957 29168
rect 63915 29119 63957 29128
rect 64011 29168 64053 29177
rect 64011 29128 64012 29168
rect 64052 29128 64053 29168
rect 64011 29119 64053 29128
rect 64107 29168 64149 29177
rect 64107 29128 64108 29168
rect 64148 29128 64149 29168
rect 64107 29119 64149 29128
rect 65643 29168 65685 29177
rect 65643 29128 65644 29168
rect 65684 29128 65685 29168
rect 65643 29119 65685 29128
rect 65835 29168 65877 29177
rect 65835 29128 65836 29168
rect 65876 29128 65877 29168
rect 65835 29119 65877 29128
rect 65923 29168 65981 29169
rect 65923 29128 65932 29168
rect 65972 29128 65981 29168
rect 65923 29127 65981 29128
rect 68035 29168 68093 29169
rect 68035 29128 68044 29168
rect 68084 29128 68093 29168
rect 68035 29127 68093 29128
rect 68899 29168 68957 29169
rect 68899 29128 68908 29168
rect 68948 29128 68957 29168
rect 68899 29127 68957 29128
rect 70347 29168 70389 29177
rect 70347 29128 70348 29168
rect 70388 29128 70389 29168
rect 70347 29119 70389 29128
rect 70443 29168 70485 29177
rect 70443 29128 70444 29168
rect 70484 29128 70485 29168
rect 70443 29119 70485 29128
rect 70539 29168 70581 29177
rect 70539 29128 70540 29168
rect 70580 29128 70581 29168
rect 73795 29168 73853 29169
rect 70539 29119 70581 29128
rect 73419 29126 73461 29135
rect 73795 29128 73804 29168
rect 73844 29128 73853 29168
rect 73795 29127 73853 29128
rect 74659 29168 74717 29169
rect 74659 29128 74668 29168
rect 74708 29128 74717 29168
rect 74659 29127 74717 29128
rect 76099 29168 76157 29169
rect 76099 29128 76108 29168
rect 76148 29128 76157 29168
rect 76099 29127 76157 29128
rect 76395 29168 76437 29177
rect 76395 29128 76396 29168
rect 76436 29128 76437 29168
rect 63339 29108 63381 29117
rect 53251 29091 53309 29092
rect 49411 29084 49469 29085
rect 49411 29044 49420 29084
rect 49460 29044 49469 29084
rect 49411 29043 49469 29044
rect 49987 29084 50045 29085
rect 49987 29044 49996 29084
rect 50036 29044 50045 29084
rect 49987 29043 50045 29044
rect 59203 29084 59261 29085
rect 59203 29044 59212 29084
rect 59252 29044 59261 29084
rect 59203 29043 59261 29044
rect 70059 29084 70101 29093
rect 73419 29086 73420 29126
rect 73460 29086 73461 29126
rect 76395 29119 76437 29128
rect 77067 29168 77109 29177
rect 77067 29128 77068 29168
rect 77108 29128 77109 29168
rect 77067 29119 77109 29128
rect 77443 29168 77501 29169
rect 77443 29128 77452 29168
rect 77492 29128 77501 29168
rect 77443 29127 77501 29128
rect 78307 29168 78365 29169
rect 78307 29128 78316 29168
rect 78356 29128 78365 29168
rect 78307 29127 78365 29128
rect 70059 29044 70060 29084
rect 70100 29044 70101 29084
rect 70059 29035 70101 29044
rect 70915 29084 70973 29085
rect 70915 29044 70924 29084
rect 70964 29044 70973 29084
rect 70915 29043 70973 29044
rect 71107 29084 71165 29085
rect 71107 29044 71116 29084
rect 71156 29044 71165 29084
rect 71107 29043 71165 29044
rect 71491 29084 71549 29085
rect 71491 29044 71500 29084
rect 71540 29044 71549 29084
rect 71491 29043 71549 29044
rect 72067 29084 72125 29085
rect 72067 29044 72076 29084
rect 72116 29044 72125 29084
rect 73419 29077 73461 29086
rect 72067 29043 72125 29044
rect 41059 29000 41117 29001
rect 41059 28960 41068 29000
rect 41108 28960 41117 29000
rect 41059 28959 41117 28960
rect 42507 29000 42549 29009
rect 42507 28960 42508 29000
rect 42548 28960 42549 29000
rect 42507 28951 42549 28960
rect 44715 29000 44757 29009
rect 44715 28960 44716 29000
rect 44756 28960 44757 29000
rect 44715 28951 44757 28960
rect 45099 29000 45141 29009
rect 45099 28960 45100 29000
rect 45140 28960 45141 29000
rect 45099 28951 45141 28960
rect 45667 29000 45725 29001
rect 45667 28960 45676 29000
rect 45716 28960 45725 29000
rect 45667 28959 45725 28960
rect 49803 29000 49845 29009
rect 49803 28960 49804 29000
rect 49844 28960 49845 29000
rect 49803 28951 49845 28960
rect 59403 29000 59445 29009
rect 59403 28960 59404 29000
rect 59444 28960 59445 29000
rect 59403 28951 59445 28960
rect 62379 29000 62421 29009
rect 62379 28960 62380 29000
rect 62420 28960 62421 29000
rect 62379 28951 62421 28960
rect 67467 29000 67509 29009
rect 67467 28960 67468 29000
rect 67508 28960 67509 29000
rect 67467 28951 67509 28960
rect 71307 29000 71349 29009
rect 71307 28960 71308 29000
rect 71348 28960 71349 29000
rect 71307 28951 71349 28960
rect 76771 29000 76829 29001
rect 76771 28960 76780 29000
rect 76820 28960 76829 29000
rect 76771 28959 76829 28960
rect 40867 28916 40925 28917
rect 40867 28876 40876 28916
rect 40916 28876 40925 28916
rect 40867 28875 40925 28876
rect 42315 28916 42357 28925
rect 42315 28876 42316 28916
rect 42356 28876 42357 28916
rect 42315 28867 42357 28876
rect 50187 28916 50229 28925
rect 50187 28876 50188 28916
rect 50228 28876 50229 28916
rect 50187 28867 50229 28876
rect 58531 28916 58589 28917
rect 58531 28876 58540 28916
rect 58580 28876 58589 28916
rect 58531 28875 58589 28876
rect 59883 28916 59925 28925
rect 59883 28876 59884 28916
rect 59924 28876 59925 28916
rect 59883 28867 59925 28876
rect 71883 28916 71925 28925
rect 71883 28876 71884 28916
rect 71924 28876 71925 28916
rect 71883 28867 71925 28876
rect 79459 28916 79517 28917
rect 79459 28876 79468 28916
rect 79508 28876 79517 28916
rect 79459 28875 79517 28876
rect 576 28748 79584 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 75112 28748
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75480 28708 79584 28748
rect 576 28684 79584 28708
rect 41067 28580 41109 28589
rect 41067 28540 41068 28580
rect 41108 28540 41109 28580
rect 41067 28531 41109 28540
rect 41643 28580 41685 28589
rect 41643 28540 41644 28580
rect 41684 28540 41685 28580
rect 41643 28531 41685 28540
rect 44619 28580 44661 28589
rect 44619 28540 44620 28580
rect 44660 28540 44661 28580
rect 44619 28531 44661 28540
rect 51339 28580 51381 28589
rect 51339 28540 51340 28580
rect 51380 28540 51381 28580
rect 51339 28531 51381 28540
rect 54603 28580 54645 28589
rect 54603 28540 54604 28580
rect 54644 28540 54645 28580
rect 54603 28531 54645 28540
rect 56035 28580 56093 28581
rect 56035 28540 56044 28580
rect 56084 28540 56093 28580
rect 56035 28539 56093 28540
rect 56235 28580 56277 28589
rect 56235 28540 56236 28580
rect 56276 28540 56277 28580
rect 56235 28531 56277 28540
rect 61035 28580 61077 28589
rect 61035 28540 61036 28580
rect 61076 28540 61077 28580
rect 61035 28531 61077 28540
rect 61611 28580 61653 28589
rect 61611 28540 61612 28580
rect 61652 28540 61653 28580
rect 61611 28531 61653 28540
rect 76779 28580 76821 28589
rect 76779 28540 76780 28580
rect 76820 28540 76821 28580
rect 76779 28531 76821 28540
rect 47595 28496 47637 28505
rect 47595 28456 47596 28496
rect 47636 28456 47637 28496
rect 47595 28447 47637 28456
rect 49323 28496 49365 28505
rect 49323 28456 49324 28496
rect 49364 28456 49365 28496
rect 49323 28447 49365 28456
rect 51723 28496 51765 28505
rect 51723 28456 51724 28496
rect 51764 28456 51765 28496
rect 51723 28447 51765 28456
rect 52299 28496 52341 28505
rect 52299 28456 52300 28496
rect 52340 28456 52341 28496
rect 52299 28447 52341 28456
rect 52491 28496 52533 28505
rect 52491 28456 52492 28496
rect 52532 28456 52533 28496
rect 52491 28447 52533 28456
rect 57771 28496 57813 28505
rect 57771 28456 57772 28496
rect 57812 28456 57813 28496
rect 57771 28447 57813 28456
rect 64483 28496 64541 28497
rect 64483 28456 64492 28496
rect 64532 28456 64541 28496
rect 64483 28455 64541 28456
rect 70915 28496 70973 28497
rect 70915 28456 70924 28496
rect 70964 28456 70973 28496
rect 70915 28455 70973 28456
rect 39523 28412 39581 28413
rect 39523 28372 39532 28412
rect 39572 28372 39581 28412
rect 39523 28371 39581 28372
rect 40099 28412 40157 28413
rect 40099 28372 40108 28412
rect 40148 28372 40157 28412
rect 40099 28371 40157 28372
rect 46243 28412 46301 28413
rect 46243 28372 46252 28412
rect 46292 28372 46301 28412
rect 46243 28371 46301 28372
rect 51139 28412 51197 28413
rect 51139 28372 51148 28412
rect 51188 28372 51197 28412
rect 51139 28371 51197 28372
rect 58915 28412 58973 28413
rect 58915 28372 58924 28412
rect 58964 28372 58973 28412
rect 58915 28371 58973 28372
rect 59587 28412 59645 28413
rect 59587 28372 59596 28412
rect 59636 28372 59645 28412
rect 59587 28371 59645 28372
rect 61219 28412 61277 28413
rect 61219 28372 61228 28412
rect 61268 28372 61277 28412
rect 61219 28371 61277 28372
rect 61411 28412 61469 28413
rect 61411 28372 61420 28412
rect 61460 28372 61469 28412
rect 61411 28371 61469 28372
rect 73803 28412 73845 28421
rect 73803 28372 73804 28412
rect 73844 28372 73845 28412
rect 73803 28363 73845 28372
rect 40299 28328 40341 28337
rect 40299 28288 40300 28328
rect 40340 28288 40341 28328
rect 40299 28279 40341 28288
rect 40491 28328 40533 28337
rect 40491 28288 40492 28328
rect 40532 28288 40533 28328
rect 40491 28279 40533 28288
rect 40579 28328 40637 28329
rect 40579 28288 40588 28328
rect 40628 28288 40637 28328
rect 40579 28287 40637 28288
rect 41067 28328 41109 28337
rect 41067 28288 41068 28328
rect 41108 28288 41109 28328
rect 41067 28279 41109 28288
rect 41259 28328 41301 28337
rect 41259 28288 41260 28328
rect 41300 28288 41301 28328
rect 41259 28279 41301 28288
rect 41347 28328 41405 28329
rect 41347 28288 41356 28328
rect 41396 28288 41405 28328
rect 41347 28287 41405 28288
rect 41547 28328 41589 28337
rect 41547 28288 41548 28328
rect 41588 28288 41589 28328
rect 41547 28279 41589 28288
rect 41731 28328 41789 28329
rect 41731 28288 41740 28328
rect 41780 28288 41789 28328
rect 41731 28287 41789 28288
rect 41931 28328 41973 28337
rect 41931 28288 41932 28328
rect 41972 28288 41973 28328
rect 41931 28279 41973 28288
rect 42307 28328 42365 28329
rect 42307 28288 42316 28328
rect 42356 28288 42365 28328
rect 42307 28287 42365 28288
rect 43212 28328 43254 28337
rect 43212 28288 43213 28328
rect 43253 28288 43254 28328
rect 43212 28279 43254 28288
rect 44619 28328 44661 28337
rect 44619 28288 44620 28328
rect 44660 28288 44661 28328
rect 44619 28279 44661 28288
rect 44811 28328 44853 28337
rect 44811 28288 44812 28328
rect 44852 28288 44853 28328
rect 44811 28279 44853 28288
rect 44899 28328 44957 28329
rect 44899 28288 44908 28328
rect 44948 28288 44957 28328
rect 44899 28287 44957 28288
rect 45099 28328 45141 28337
rect 45099 28288 45100 28328
rect 45140 28288 45141 28328
rect 45099 28279 45141 28288
rect 45195 28328 45237 28337
rect 45195 28288 45196 28328
rect 45236 28288 45237 28328
rect 45195 28279 45237 28288
rect 45291 28328 45333 28337
rect 45291 28288 45292 28328
rect 45332 28288 45333 28328
rect 45291 28279 45333 28288
rect 45387 28328 45429 28337
rect 45387 28288 45388 28328
rect 45428 28288 45429 28328
rect 45387 28279 45429 28288
rect 45579 28328 45621 28337
rect 45579 28288 45580 28328
rect 45620 28288 45621 28328
rect 45579 28279 45621 28288
rect 45771 28328 45813 28337
rect 45771 28288 45772 28328
rect 45812 28288 45813 28328
rect 45771 28279 45813 28288
rect 45859 28328 45917 28329
rect 45859 28288 45868 28328
rect 45908 28288 45917 28328
rect 45859 28287 45917 28288
rect 46627 28328 46685 28329
rect 46627 28288 46636 28328
rect 46676 28288 46685 28328
rect 46627 28287 46685 28288
rect 46827 28328 46869 28337
rect 46827 28288 46828 28328
rect 46868 28288 46869 28328
rect 46827 28279 46869 28288
rect 49995 28328 50037 28337
rect 49995 28288 49996 28328
rect 50036 28288 50037 28328
rect 49995 28279 50037 28288
rect 50187 28328 50229 28337
rect 50187 28288 50188 28328
rect 50228 28288 50229 28328
rect 50187 28279 50229 28288
rect 50275 28328 50333 28329
rect 50275 28288 50284 28328
rect 50324 28288 50333 28328
rect 50275 28287 50333 28288
rect 50475 28328 50517 28337
rect 50475 28288 50476 28328
rect 50516 28288 50517 28328
rect 50475 28279 50517 28288
rect 50571 28328 50613 28337
rect 50571 28288 50572 28328
rect 50612 28288 50613 28328
rect 50571 28279 50613 28288
rect 50667 28328 50709 28337
rect 50667 28288 50668 28328
rect 50708 28288 50709 28328
rect 50667 28279 50709 28288
rect 50763 28328 50805 28337
rect 50763 28288 50764 28328
rect 50804 28288 50805 28328
rect 50763 28279 50805 28288
rect 51619 28328 51677 28329
rect 51619 28288 51628 28328
rect 51668 28288 51677 28328
rect 51619 28287 51677 28288
rect 51819 28328 51861 28337
rect 51819 28288 51820 28328
rect 51860 28288 51861 28328
rect 51819 28279 51861 28288
rect 52963 28328 53021 28329
rect 52963 28288 52972 28328
rect 53012 28288 53021 28328
rect 52963 28287 53021 28288
rect 55363 28328 55421 28329
rect 55363 28288 55372 28328
rect 55412 28288 55421 28328
rect 55363 28287 55421 28288
rect 55659 28328 55701 28337
rect 55659 28288 55660 28328
rect 55700 28288 55701 28328
rect 55659 28279 55701 28288
rect 55755 28328 55797 28337
rect 55755 28288 55756 28328
rect 55796 28288 55797 28328
rect 55755 28279 55797 28288
rect 56235 28328 56277 28337
rect 56235 28288 56236 28328
rect 56276 28288 56277 28328
rect 56235 28279 56277 28288
rect 56427 28328 56469 28337
rect 56427 28288 56428 28328
rect 56468 28288 56469 28328
rect 56427 28279 56469 28288
rect 56515 28328 56573 28329
rect 56515 28288 56524 28328
rect 56564 28288 56573 28328
rect 56515 28287 56573 28288
rect 56707 28328 56765 28329
rect 56707 28288 56716 28328
rect 56756 28288 56765 28328
rect 56707 28287 56765 28288
rect 56907 28328 56949 28337
rect 56907 28288 56908 28328
rect 56948 28288 56949 28328
rect 56907 28279 56949 28288
rect 59115 28328 59157 28337
rect 59115 28288 59116 28328
rect 59156 28288 59157 28328
rect 59115 28279 59157 28288
rect 59211 28328 59253 28337
rect 59211 28288 59212 28328
rect 59252 28288 59253 28328
rect 59211 28279 59253 28288
rect 59307 28328 59349 28337
rect 59307 28288 59308 28328
rect 59348 28288 59349 28328
rect 59307 28279 59349 28288
rect 60171 28328 60213 28337
rect 60171 28288 60172 28328
rect 60212 28288 60213 28328
rect 60171 28279 60213 28288
rect 60363 28328 60405 28337
rect 60363 28288 60364 28328
rect 60404 28288 60405 28328
rect 60363 28279 60405 28288
rect 60451 28328 60509 28329
rect 60451 28288 60460 28328
rect 60500 28288 60509 28328
rect 60451 28287 60509 28288
rect 60651 28328 60693 28337
rect 60651 28288 60652 28328
rect 60692 28288 60693 28328
rect 60651 28279 60693 28288
rect 60747 28328 60789 28337
rect 60747 28288 60748 28328
rect 60788 28288 60789 28328
rect 60747 28279 60789 28288
rect 60835 28328 60893 28329
rect 60835 28288 60844 28328
rect 60884 28288 60893 28328
rect 60835 28287 60893 28288
rect 62275 28328 62333 28329
rect 62275 28288 62284 28328
rect 62324 28288 62333 28328
rect 62275 28287 62333 28288
rect 63139 28328 63197 28329
rect 63139 28288 63148 28328
rect 63188 28288 63197 28328
rect 63139 28287 63197 28288
rect 64779 28328 64821 28337
rect 64779 28288 64780 28328
rect 64820 28288 64821 28328
rect 64779 28279 64821 28288
rect 64875 28328 64917 28337
rect 64875 28288 64876 28328
rect 64916 28288 64917 28328
rect 64875 28279 64917 28288
rect 65155 28328 65213 28329
rect 65155 28288 65164 28328
rect 65204 28288 65213 28328
rect 65155 28287 65213 28288
rect 66115 28328 66173 28329
rect 66115 28288 66124 28328
rect 66164 28288 66173 28328
rect 66115 28287 66173 28288
rect 66979 28328 67037 28329
rect 66979 28288 66988 28328
rect 67028 28288 67037 28328
rect 66979 28287 67037 28288
rect 70243 28328 70301 28329
rect 70243 28288 70252 28328
rect 70292 28288 70301 28328
rect 70243 28287 70301 28288
rect 70539 28328 70581 28337
rect 70539 28288 70540 28328
rect 70580 28288 70581 28328
rect 70539 28279 70581 28288
rect 70635 28328 70677 28337
rect 70635 28288 70636 28328
rect 70676 28288 70677 28328
rect 70635 28279 70677 28288
rect 71779 28328 71837 28329
rect 71779 28288 71788 28328
rect 71828 28288 71837 28328
rect 71779 28287 71837 28288
rect 72643 28328 72701 28329
rect 72643 28288 72652 28328
rect 72692 28288 72701 28328
rect 72643 28287 72701 28288
rect 75243 28328 75285 28337
rect 75243 28288 75244 28328
rect 75284 28288 75285 28328
rect 75243 28279 75285 28288
rect 75435 28328 75477 28337
rect 75435 28288 75436 28328
rect 75476 28288 75477 28328
rect 75435 28279 75477 28288
rect 75523 28328 75581 28329
rect 75523 28288 75532 28328
rect 75572 28288 75581 28328
rect 75523 28287 75581 28288
rect 76779 28328 76821 28337
rect 76779 28288 76780 28328
rect 76820 28288 76821 28328
rect 76779 28279 76821 28288
rect 76971 28328 77013 28337
rect 76971 28288 76972 28328
rect 77012 28288 77013 28328
rect 76971 28279 77013 28288
rect 77059 28328 77117 28329
rect 77059 28288 77068 28328
rect 77108 28288 77117 28328
rect 77059 28287 77117 28288
rect 77251 28328 77309 28329
rect 77251 28288 77260 28328
rect 77300 28288 77309 28328
rect 77251 28287 77309 28288
rect 77451 28328 77493 28337
rect 77451 28288 77452 28328
rect 77492 28288 77493 28328
rect 77451 28279 77493 28288
rect 46731 28244 46773 28253
rect 46731 28204 46732 28244
rect 46772 28204 46773 28244
rect 46731 28195 46773 28204
rect 56811 28244 56853 28253
rect 56811 28204 56812 28244
rect 56852 28204 56853 28244
rect 56811 28195 56853 28204
rect 61899 28244 61941 28253
rect 61899 28204 61900 28244
rect 61940 28204 61941 28244
rect 61899 28195 61941 28204
rect 65739 28244 65781 28253
rect 65739 28204 65740 28244
rect 65780 28204 65781 28244
rect 65739 28195 65781 28204
rect 71403 28244 71445 28253
rect 71403 28204 71404 28244
rect 71444 28204 71445 28244
rect 71403 28195 71445 28204
rect 75339 28244 75381 28253
rect 75339 28204 75340 28244
rect 75380 28204 75381 28244
rect 75339 28195 75381 28204
rect 77355 28244 77397 28253
rect 77355 28204 77356 28244
rect 77396 28204 77397 28244
rect 77355 28195 77397 28204
rect 39723 28160 39765 28169
rect 39723 28120 39724 28160
rect 39764 28120 39765 28160
rect 39723 28111 39765 28120
rect 39915 28160 39957 28169
rect 39915 28120 39916 28160
rect 39956 28120 39957 28160
rect 39915 28111 39957 28120
rect 40387 28160 40445 28161
rect 40387 28120 40396 28160
rect 40436 28120 40445 28160
rect 40387 28119 40445 28120
rect 44323 28160 44381 28161
rect 44323 28120 44332 28160
rect 44372 28120 44381 28160
rect 44323 28119 44381 28120
rect 45667 28160 45725 28161
rect 45667 28120 45676 28160
rect 45716 28120 45725 28160
rect 45667 28119 45725 28120
rect 46059 28160 46101 28169
rect 46059 28120 46060 28160
rect 46100 28120 46101 28160
rect 46059 28111 46101 28120
rect 50083 28160 50141 28161
rect 50083 28120 50092 28160
rect 50132 28120 50141 28160
rect 50083 28119 50141 28120
rect 58731 28160 58773 28169
rect 58731 28120 58732 28160
rect 58772 28120 58773 28160
rect 58731 28111 58773 28120
rect 59395 28160 59453 28161
rect 59395 28120 59404 28160
rect 59444 28120 59453 28160
rect 59395 28119 59453 28120
rect 59787 28160 59829 28169
rect 59787 28120 59788 28160
rect 59828 28120 59829 28160
rect 59787 28111 59829 28120
rect 60259 28160 60317 28161
rect 60259 28120 60268 28160
rect 60308 28120 60317 28160
rect 60259 28119 60317 28120
rect 61035 28160 61077 28169
rect 61035 28120 61036 28160
rect 61076 28120 61077 28160
rect 61035 28111 61077 28120
rect 64291 28160 64349 28161
rect 64291 28120 64300 28160
rect 64340 28120 64349 28160
rect 64291 28119 64349 28120
rect 68131 28160 68189 28161
rect 68131 28120 68140 28160
rect 68180 28120 68189 28160
rect 68131 28119 68189 28120
rect 576 27992 79584 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 76352 27992
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76720 27952 79584 27992
rect 576 27928 79584 27952
rect 3819 27824 3861 27833
rect 3819 27784 3820 27824
rect 3860 27784 3861 27824
rect 3819 27775 3861 27784
rect 41451 27824 41493 27833
rect 41451 27784 41452 27824
rect 41492 27784 41493 27824
rect 41451 27775 41493 27784
rect 43555 27824 43613 27825
rect 43555 27784 43564 27824
rect 43604 27784 43613 27824
rect 43555 27783 43613 27784
rect 51235 27824 51293 27825
rect 51235 27784 51244 27824
rect 51284 27784 51293 27824
rect 51235 27783 51293 27784
rect 59683 27824 59741 27825
rect 59683 27784 59692 27824
rect 59732 27784 59741 27824
rect 59683 27783 59741 27784
rect 63907 27824 63965 27825
rect 63907 27784 63916 27824
rect 63956 27784 63965 27824
rect 63907 27783 63965 27784
rect 71107 27824 71165 27825
rect 71107 27784 71116 27824
rect 71156 27784 71165 27824
rect 71107 27783 71165 27784
rect 37803 27740 37845 27749
rect 37803 27700 37804 27740
rect 37844 27700 37845 27740
rect 37803 27691 37845 27700
rect 40491 27740 40533 27749
rect 40491 27700 40492 27740
rect 40532 27700 40533 27740
rect 40491 27691 40533 27700
rect 45963 27740 46005 27749
rect 45963 27700 45964 27740
rect 46004 27700 46005 27740
rect 45963 27691 46005 27700
rect 46635 27740 46677 27749
rect 46635 27700 46636 27740
rect 46676 27700 46677 27740
rect 46635 27691 46677 27700
rect 47691 27740 47733 27749
rect 47691 27700 47692 27740
rect 47732 27700 47733 27740
rect 47691 27691 47733 27700
rect 48843 27740 48885 27749
rect 48843 27700 48844 27740
rect 48884 27700 48885 27740
rect 48843 27691 48885 27700
rect 51627 27740 51669 27749
rect 51627 27700 51628 27740
rect 51668 27700 51669 27740
rect 51627 27691 51669 27700
rect 52011 27740 52053 27749
rect 52011 27700 52012 27740
rect 52052 27700 52053 27740
rect 52011 27691 52053 27700
rect 57291 27740 57333 27749
rect 57291 27700 57292 27740
rect 57332 27700 57333 27740
rect 57291 27691 57333 27700
rect 59979 27740 60021 27749
rect 59979 27700 59980 27740
rect 60020 27700 60021 27740
rect 59979 27691 60021 27700
rect 60555 27740 60597 27749
rect 60555 27700 60556 27740
rect 60596 27700 60597 27740
rect 60555 27691 60597 27700
rect 70731 27740 70773 27749
rect 70731 27700 70732 27740
rect 70772 27700 70773 27740
rect 70731 27691 70773 27700
rect 71691 27669 71733 27678
rect 3715 27656 3773 27657
rect 3715 27616 3724 27656
rect 3764 27616 3773 27656
rect 3715 27615 3773 27616
rect 38179 27656 38237 27657
rect 38179 27616 38188 27656
rect 38228 27616 38237 27656
rect 38179 27615 38237 27616
rect 39043 27656 39101 27657
rect 39043 27616 39052 27656
rect 39092 27616 39101 27656
rect 39043 27615 39101 27616
rect 40395 27656 40437 27665
rect 40395 27616 40396 27656
rect 40436 27616 40437 27656
rect 40395 27607 40437 27616
rect 40587 27656 40629 27665
rect 40587 27616 40588 27656
rect 40628 27616 40629 27656
rect 40587 27607 40629 27616
rect 40675 27656 40733 27657
rect 40675 27616 40684 27656
rect 40724 27616 40733 27656
rect 40675 27615 40733 27616
rect 41059 27656 41117 27657
rect 41059 27616 41068 27656
rect 41108 27616 41117 27656
rect 41059 27615 41117 27616
rect 41259 27656 41301 27665
rect 41259 27616 41260 27656
rect 41300 27616 41301 27656
rect 41259 27607 41301 27616
rect 44707 27656 44765 27657
rect 44707 27616 44716 27656
rect 44756 27616 44765 27656
rect 44707 27615 44765 27616
rect 45571 27656 45629 27657
rect 45571 27616 45580 27656
rect 45620 27616 45629 27656
rect 45571 27615 45629 27616
rect 46243 27656 46301 27657
rect 46243 27616 46252 27656
rect 46292 27616 46301 27656
rect 46243 27615 46301 27616
rect 46539 27656 46581 27665
rect 46539 27616 46540 27656
rect 46580 27616 46581 27656
rect 46539 27607 46581 27616
rect 47115 27656 47157 27665
rect 47115 27616 47116 27656
rect 47156 27616 47157 27656
rect 47115 27607 47157 27616
rect 47307 27656 47349 27665
rect 47307 27616 47308 27656
rect 47348 27616 47349 27656
rect 47307 27607 47349 27616
rect 47395 27656 47453 27657
rect 47395 27616 47404 27656
rect 47444 27616 47453 27656
rect 47395 27615 47453 27616
rect 47587 27656 47645 27657
rect 47587 27616 47596 27656
rect 47636 27616 47645 27656
rect 47587 27615 47645 27616
rect 47787 27656 47829 27665
rect 47787 27616 47788 27656
rect 47828 27616 47829 27656
rect 47787 27607 47829 27616
rect 47971 27656 48029 27657
rect 47971 27616 47980 27656
rect 48020 27616 48029 27656
rect 47971 27615 48029 27616
rect 49219 27656 49277 27657
rect 49219 27616 49228 27656
rect 49268 27616 49277 27656
rect 49219 27615 49277 27616
rect 50083 27656 50141 27657
rect 50083 27616 50092 27656
rect 50132 27616 50141 27656
rect 50083 27615 50141 27616
rect 51531 27656 51573 27665
rect 51531 27616 51532 27656
rect 51572 27616 51573 27656
rect 51531 27607 51573 27616
rect 51723 27656 51765 27665
rect 51723 27616 51724 27656
rect 51764 27616 51765 27656
rect 51723 27607 51765 27616
rect 51811 27656 51869 27657
rect 51811 27616 51820 27656
rect 51860 27616 51869 27656
rect 51811 27615 51869 27616
rect 52387 27656 52445 27657
rect 52387 27616 52396 27656
rect 52436 27616 52445 27656
rect 52387 27615 52445 27616
rect 53292 27656 53334 27665
rect 53292 27616 53293 27656
rect 53333 27616 53334 27656
rect 53292 27607 53334 27616
rect 54603 27656 54645 27665
rect 54603 27616 54604 27656
rect 54644 27616 54645 27656
rect 54603 27607 54645 27616
rect 54795 27656 54837 27665
rect 54795 27616 54796 27656
rect 54836 27616 54837 27656
rect 54795 27607 54837 27616
rect 54883 27656 54941 27657
rect 54883 27616 54892 27656
rect 54932 27616 54941 27656
rect 54883 27615 54941 27616
rect 55179 27656 55221 27665
rect 55179 27616 55180 27656
rect 55220 27616 55221 27656
rect 55179 27607 55221 27616
rect 55371 27656 55413 27665
rect 55371 27616 55372 27656
rect 55412 27616 55413 27656
rect 55371 27607 55413 27616
rect 55459 27656 55517 27657
rect 55459 27616 55468 27656
rect 55508 27616 55517 27656
rect 55459 27615 55517 27616
rect 55659 27656 55701 27665
rect 55659 27616 55660 27656
rect 55700 27616 55701 27656
rect 55659 27607 55701 27616
rect 55755 27656 55797 27665
rect 55755 27616 55756 27656
rect 55796 27616 55797 27656
rect 55755 27607 55797 27616
rect 55851 27656 55893 27665
rect 55851 27616 55852 27656
rect 55892 27616 55893 27656
rect 55851 27607 55893 27616
rect 55947 27656 55989 27665
rect 55947 27616 55948 27656
rect 55988 27616 55989 27656
rect 55947 27607 55989 27616
rect 57667 27656 57725 27657
rect 57667 27616 57676 27656
rect 57716 27616 57725 27656
rect 57667 27615 57725 27616
rect 58531 27656 58589 27657
rect 58531 27616 58540 27656
rect 58580 27616 58589 27656
rect 58531 27615 58589 27616
rect 59883 27656 59925 27665
rect 59883 27616 59884 27656
rect 59924 27616 59925 27656
rect 59883 27607 59925 27616
rect 60075 27656 60117 27665
rect 60075 27616 60076 27656
rect 60116 27616 60117 27656
rect 60075 27607 60117 27616
rect 60163 27656 60221 27657
rect 60163 27616 60172 27656
rect 60212 27616 60221 27656
rect 60163 27615 60221 27616
rect 60931 27656 60989 27657
rect 60931 27616 60940 27656
rect 60980 27616 60989 27656
rect 60931 27615 60989 27616
rect 61795 27656 61853 27657
rect 61795 27616 61804 27656
rect 61844 27616 61853 27656
rect 61795 27615 61853 27616
rect 63715 27656 63773 27657
rect 63715 27616 63724 27656
rect 63764 27616 63773 27656
rect 63715 27615 63773 27616
rect 63819 27656 63861 27665
rect 63819 27616 63820 27656
rect 63860 27616 63861 27656
rect 63819 27607 63861 27616
rect 64011 27656 64053 27665
rect 64011 27616 64012 27656
rect 64052 27616 64053 27656
rect 64011 27607 64053 27616
rect 64779 27656 64821 27665
rect 64779 27616 64780 27656
rect 64820 27616 64821 27656
rect 64779 27607 64821 27616
rect 64875 27656 64917 27665
rect 64875 27616 64876 27656
rect 64916 27616 64917 27656
rect 64875 27607 64917 27616
rect 64963 27656 65021 27657
rect 64963 27616 64972 27656
rect 65012 27616 65021 27656
rect 64963 27615 65021 27616
rect 65163 27656 65205 27665
rect 65163 27616 65164 27656
rect 65204 27616 65205 27656
rect 65163 27607 65205 27616
rect 65355 27656 65397 27665
rect 65355 27616 65356 27656
rect 65396 27616 65397 27656
rect 65355 27607 65397 27616
rect 65443 27656 65501 27657
rect 65443 27616 65452 27656
rect 65492 27616 65501 27656
rect 65443 27615 65501 27616
rect 65635 27656 65693 27657
rect 65635 27616 65644 27656
rect 65684 27616 65693 27656
rect 65635 27615 65693 27616
rect 65835 27656 65877 27665
rect 65835 27616 65836 27656
rect 65876 27616 65877 27656
rect 65835 27607 65877 27616
rect 69579 27656 69621 27665
rect 69579 27616 69580 27656
rect 69620 27616 69621 27656
rect 69579 27607 69621 27616
rect 69771 27656 69813 27665
rect 69771 27616 69772 27656
rect 69812 27616 69813 27656
rect 69771 27607 69813 27616
rect 69859 27656 69917 27657
rect 69859 27616 69868 27656
rect 69908 27616 69917 27656
rect 69859 27615 69917 27616
rect 70059 27656 70101 27665
rect 70059 27616 70060 27656
rect 70100 27616 70101 27656
rect 70059 27607 70101 27616
rect 70251 27656 70293 27665
rect 70251 27616 70252 27656
rect 70292 27616 70293 27656
rect 70251 27607 70293 27616
rect 70339 27656 70397 27657
rect 70339 27616 70348 27656
rect 70388 27616 70397 27656
rect 70339 27615 70397 27616
rect 70627 27656 70685 27657
rect 70627 27616 70636 27656
rect 70676 27616 70685 27656
rect 70627 27615 70685 27616
rect 70827 27656 70869 27665
rect 70827 27616 70828 27656
rect 70868 27616 70869 27656
rect 70827 27607 70869 27616
rect 71019 27656 71061 27665
rect 71019 27616 71020 27656
rect 71060 27616 71061 27656
rect 71019 27607 71061 27616
rect 71211 27656 71253 27665
rect 71211 27616 71212 27656
rect 71252 27616 71253 27656
rect 71211 27607 71253 27616
rect 71299 27656 71357 27657
rect 71299 27616 71308 27656
rect 71348 27616 71357 27656
rect 71299 27615 71357 27616
rect 71491 27656 71549 27657
rect 71491 27616 71500 27656
rect 71540 27616 71549 27656
rect 71691 27629 71692 27669
rect 71732 27629 71733 27669
rect 71691 27620 71733 27629
rect 74859 27656 74901 27665
rect 71491 27615 71549 27616
rect 74859 27616 74860 27656
rect 74900 27616 74901 27656
rect 74859 27607 74901 27616
rect 75051 27656 75093 27665
rect 75051 27616 75052 27656
rect 75092 27616 75093 27656
rect 75051 27607 75093 27616
rect 75139 27656 75197 27657
rect 75139 27616 75148 27656
rect 75188 27616 75197 27656
rect 75139 27615 75197 27616
rect 75435 27656 75477 27665
rect 75435 27616 75436 27656
rect 75476 27616 75477 27656
rect 75435 27607 75477 27616
rect 75627 27656 75669 27665
rect 75627 27616 75628 27656
rect 75668 27616 75669 27656
rect 75627 27607 75669 27616
rect 75715 27656 75773 27657
rect 75715 27616 75724 27656
rect 75764 27616 75773 27656
rect 75715 27615 75773 27616
rect 76675 27656 76733 27657
rect 76675 27616 76684 27656
rect 76724 27616 76733 27656
rect 76675 27615 76733 27616
rect 76779 27656 76821 27665
rect 76779 27616 76780 27656
rect 76820 27616 76821 27656
rect 76779 27607 76821 27616
rect 76875 27656 76917 27665
rect 76875 27616 76876 27656
rect 76916 27616 76917 27656
rect 76875 27607 76917 27616
rect 77155 27656 77213 27657
rect 77155 27616 77164 27656
rect 77204 27616 77213 27656
rect 77155 27615 77213 27616
rect 77355 27656 77397 27665
rect 77355 27616 77356 27656
rect 77396 27616 77397 27656
rect 77355 27607 77397 27616
rect 41635 27572 41693 27573
rect 41635 27532 41644 27572
rect 41684 27532 41693 27572
rect 41635 27531 41693 27532
rect 65739 27572 65781 27581
rect 65739 27532 65740 27572
rect 65780 27532 65781 27572
rect 65739 27523 65781 27532
rect 67555 27572 67613 27573
rect 67555 27532 67564 27572
rect 67604 27532 67613 27572
rect 67555 27531 67613 27532
rect 46915 27488 46973 27489
rect 46915 27448 46924 27488
rect 46964 27448 46973 27488
rect 46915 27447 46973 27448
rect 54603 27488 54645 27497
rect 54603 27448 54604 27488
rect 54644 27448 54645 27488
rect 54603 27439 54645 27448
rect 56139 27488 56181 27497
rect 56139 27448 56140 27488
rect 56180 27448 56181 27488
rect 56139 27439 56181 27448
rect 59683 27488 59741 27489
rect 59683 27448 59692 27488
rect 59732 27448 59741 27488
rect 59683 27447 59741 27448
rect 65163 27488 65205 27497
rect 65163 27448 65164 27488
rect 65204 27448 65205 27488
rect 65163 27439 65205 27448
rect 66219 27488 66261 27497
rect 66219 27448 66220 27488
rect 66260 27448 66261 27488
rect 66219 27439 66261 27448
rect 69387 27488 69429 27497
rect 69387 27448 69388 27488
rect 69428 27448 69429 27488
rect 69387 27439 69429 27448
rect 69579 27488 69621 27497
rect 69579 27448 69580 27488
rect 69620 27448 69621 27488
rect 69579 27439 69621 27448
rect 70059 27488 70101 27497
rect 70059 27448 70060 27488
rect 70100 27448 70101 27488
rect 70059 27439 70101 27448
rect 71883 27488 71925 27497
rect 71883 27448 71884 27488
rect 71924 27448 71925 27488
rect 71883 27439 71925 27448
rect 73515 27488 73557 27497
rect 73515 27448 73516 27488
rect 73556 27448 73557 27488
rect 73515 27439 73557 27448
rect 77547 27488 77589 27497
rect 77547 27448 77548 27488
rect 77588 27448 77589 27488
rect 77547 27439 77589 27448
rect 3819 27404 3861 27413
rect 3819 27364 3820 27404
rect 3860 27364 3861 27404
rect 3819 27355 3861 27364
rect 40195 27404 40253 27405
rect 40195 27364 40204 27404
rect 40244 27364 40253 27404
rect 40195 27363 40253 27364
rect 41163 27404 41205 27413
rect 41163 27364 41164 27404
rect 41204 27364 41205 27404
rect 41163 27355 41205 27364
rect 41451 27404 41493 27413
rect 41451 27364 41452 27404
rect 41492 27364 41493 27404
rect 41451 27355 41493 27364
rect 47115 27404 47157 27413
rect 47115 27364 47116 27404
rect 47156 27364 47157 27404
rect 47115 27355 47157 27364
rect 51235 27404 51293 27405
rect 51235 27364 51244 27404
rect 51284 27364 51293 27404
rect 51235 27363 51293 27364
rect 54403 27404 54461 27405
rect 54403 27364 54412 27404
rect 54452 27364 54461 27404
rect 54403 27363 54461 27364
rect 55179 27404 55221 27413
rect 55179 27364 55180 27404
rect 55220 27364 55221 27404
rect 55179 27355 55221 27364
rect 62947 27404 63005 27405
rect 62947 27364 62956 27404
rect 62996 27364 63005 27404
rect 62947 27363 63005 27364
rect 67371 27404 67413 27413
rect 67371 27364 67372 27404
rect 67412 27364 67413 27404
rect 67371 27355 67413 27364
rect 71595 27404 71637 27413
rect 71595 27364 71596 27404
rect 71636 27364 71637 27404
rect 71595 27355 71637 27364
rect 74859 27404 74901 27413
rect 74859 27364 74860 27404
rect 74900 27364 74901 27404
rect 74859 27355 74901 27364
rect 75435 27404 75477 27413
rect 75435 27364 75436 27404
rect 75476 27364 75477 27404
rect 75435 27355 75477 27364
rect 77259 27404 77301 27413
rect 77259 27364 77260 27404
rect 77300 27364 77301 27404
rect 77259 27355 77301 27364
rect 576 27236 79584 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 75112 27236
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75480 27196 79584 27236
rect 576 27172 79584 27196
rect 39723 27068 39765 27077
rect 39723 27028 39724 27068
rect 39764 27028 39765 27068
rect 39723 27019 39765 27028
rect 41155 27068 41213 27069
rect 41155 27028 41164 27068
rect 41204 27028 41213 27068
rect 41155 27027 41213 27028
rect 49507 27068 49565 27069
rect 49507 27028 49516 27068
rect 49556 27028 49565 27068
rect 49507 27027 49565 27028
rect 51811 27068 51869 27069
rect 51811 27028 51820 27068
rect 51860 27028 51869 27068
rect 51811 27027 51869 27028
rect 52107 27068 52149 27077
rect 52107 27028 52108 27068
rect 52148 27028 52149 27068
rect 52107 27019 52149 27028
rect 54211 27068 54269 27069
rect 54211 27028 54220 27068
rect 54260 27028 54269 27068
rect 54211 27027 54269 27028
rect 58539 27068 58581 27077
rect 58539 27028 58540 27068
rect 58580 27028 58581 27068
rect 58539 27019 58581 27028
rect 60163 27068 60221 27069
rect 60163 27028 60172 27068
rect 60212 27028 60221 27068
rect 60163 27027 60221 27028
rect 60843 27068 60885 27077
rect 60843 27028 60844 27068
rect 60884 27028 60885 27068
rect 60843 27019 60885 27028
rect 63819 27068 63861 27077
rect 63819 27028 63820 27068
rect 63860 27028 63861 27068
rect 63819 27019 63861 27028
rect 68811 27068 68853 27077
rect 68811 27028 68812 27068
rect 68852 27028 68853 27068
rect 68811 27019 68853 27028
rect 71979 27068 72021 27077
rect 71979 27028 71980 27068
rect 72020 27028 72021 27068
rect 71979 27019 72021 27028
rect 72171 27068 72213 27077
rect 72171 27028 72172 27068
rect 72212 27028 72213 27068
rect 72171 27019 72213 27028
rect 76867 27068 76925 27069
rect 76867 27028 76876 27068
rect 76916 27028 76925 27068
rect 76867 27027 76925 27028
rect 35115 26984 35157 26993
rect 35115 26944 35116 26984
rect 35156 26944 35157 26984
rect 35115 26935 35157 26944
rect 38283 26984 38325 26993
rect 38283 26944 38284 26984
rect 38324 26944 38325 26984
rect 38283 26935 38325 26944
rect 39339 26984 39381 26993
rect 39339 26944 39340 26984
rect 39380 26944 39381 26984
rect 39339 26935 39381 26944
rect 58155 26984 58197 26993
rect 58155 26944 58156 26984
rect 58196 26944 58197 26984
rect 58155 26935 58197 26944
rect 61131 26984 61173 26993
rect 61131 26944 61132 26984
rect 61172 26944 61173 26984
rect 61131 26935 61173 26944
rect 62091 26984 62133 26993
rect 62091 26944 62092 26984
rect 62132 26944 62133 26984
rect 62091 26935 62133 26944
rect 50397 26903 50439 26912
rect 39139 26900 39197 26901
rect 39139 26860 39148 26900
rect 39188 26860 39197 26900
rect 39139 26859 39197 26860
rect 39523 26900 39581 26901
rect 39523 26860 39532 26900
rect 39572 26860 39581 26900
rect 39523 26859 39581 26860
rect 50397 26863 50398 26903
rect 50438 26863 50439 26903
rect 50397 26854 50439 26863
rect 57955 26900 58013 26901
rect 57955 26860 57964 26900
rect 58004 26860 58013 26900
rect 57955 26859 58013 26860
rect 58339 26900 58397 26901
rect 58339 26860 58348 26900
rect 58388 26860 58397 26900
rect 58339 26859 58397 26860
rect 60355 26900 60413 26901
rect 60355 26860 60364 26900
rect 60404 26860 60413 26900
rect 60355 26859 60413 26860
rect 68995 26900 69053 26901
rect 68995 26860 69004 26900
rect 69044 26860 69053 26900
rect 68995 26859 69053 26860
rect 71779 26900 71837 26901
rect 71779 26860 71788 26900
rect 71828 26860 71837 26900
rect 71779 26859 71837 26860
rect 72355 26900 72413 26901
rect 72355 26860 72364 26900
rect 72404 26860 72413 26900
rect 72355 26859 72413 26860
rect 75435 26900 75477 26909
rect 75435 26860 75436 26900
rect 75476 26860 75477 26900
rect 73411 26852 73469 26853
rect 50571 26827 50613 26836
rect 35011 26816 35069 26817
rect 35011 26776 35020 26816
rect 35060 26776 35069 26816
rect 35011 26775 35069 26776
rect 35211 26816 35253 26825
rect 35211 26776 35212 26816
rect 35252 26776 35253 26816
rect 35211 26767 35253 26776
rect 36067 26816 36125 26817
rect 36067 26776 36076 26816
rect 36116 26776 36125 26816
rect 36067 26775 36125 26776
rect 36931 26816 36989 26817
rect 36931 26776 36940 26816
rect 36980 26776 36989 26816
rect 36931 26775 36989 26776
rect 39915 26816 39957 26825
rect 39915 26776 39916 26816
rect 39956 26776 39957 26816
rect 39915 26767 39957 26776
rect 40011 26816 40053 26825
rect 40011 26776 40012 26816
rect 40052 26776 40053 26816
rect 40011 26767 40053 26776
rect 40107 26816 40149 26825
rect 40107 26776 40108 26816
rect 40148 26776 40149 26816
rect 40107 26767 40149 26776
rect 40203 26816 40245 26825
rect 40203 26776 40204 26816
rect 40244 26776 40245 26816
rect 40203 26767 40245 26776
rect 40483 26816 40541 26817
rect 40483 26776 40492 26816
rect 40532 26776 40541 26816
rect 40483 26775 40541 26776
rect 40779 26816 40821 26825
rect 40779 26776 40780 26816
rect 40820 26776 40821 26816
rect 40779 26767 40821 26776
rect 40875 26816 40917 26825
rect 40875 26776 40876 26816
rect 40916 26776 40917 26816
rect 40875 26767 40917 26776
rect 41347 26816 41405 26817
rect 41347 26776 41356 26816
rect 41396 26776 41405 26816
rect 41347 26775 41405 26776
rect 41547 26816 41589 26825
rect 41547 26776 41548 26816
rect 41588 26776 41589 26816
rect 41547 26767 41589 26776
rect 42115 26816 42173 26817
rect 42115 26776 42124 26816
rect 42164 26776 42173 26816
rect 42115 26775 42173 26776
rect 42979 26816 43037 26817
rect 42979 26776 42988 26816
rect 43028 26776 43037 26816
rect 42979 26775 43037 26776
rect 45387 26816 45429 26825
rect 45387 26776 45388 26816
rect 45428 26776 45429 26816
rect 45387 26767 45429 26776
rect 46819 26816 46877 26817
rect 46819 26776 46828 26816
rect 46868 26776 46877 26816
rect 46819 26775 46877 26776
rect 47115 26816 47157 26825
rect 47115 26776 47116 26816
rect 47156 26776 47157 26816
rect 47115 26767 47157 26776
rect 47491 26816 47549 26817
rect 47491 26776 47500 26816
rect 47540 26776 47549 26816
rect 47491 26775 47549 26776
rect 48355 26816 48413 26817
rect 48355 26776 48364 26816
rect 48404 26776 48413 26816
rect 50571 26787 50572 26827
rect 50612 26787 50613 26827
rect 50571 26778 50613 26787
rect 50763 26816 50805 26825
rect 48355 26775 48413 26776
rect 50763 26776 50764 26816
rect 50804 26776 50805 26816
rect 50763 26767 50805 26776
rect 50851 26816 50909 26817
rect 50851 26776 50860 26816
rect 50900 26776 50909 26816
rect 50851 26775 50909 26776
rect 51139 26816 51197 26817
rect 51139 26776 51148 26816
rect 51188 26776 51197 26816
rect 51139 26775 51197 26776
rect 51435 26816 51477 26825
rect 51435 26776 51436 26816
rect 51476 26776 51477 26816
rect 51435 26767 51477 26776
rect 51531 26816 51573 26825
rect 51531 26776 51532 26816
rect 51572 26776 51573 26816
rect 51531 26767 51573 26776
rect 52003 26816 52061 26817
rect 52003 26776 52012 26816
rect 52052 26776 52061 26816
rect 52003 26775 52061 26776
rect 52203 26816 52245 26825
rect 52203 26776 52204 26816
rect 52244 26776 52245 26816
rect 52203 26767 52245 26776
rect 55363 26816 55421 26817
rect 55363 26776 55372 26816
rect 55412 26776 55421 26816
rect 55363 26775 55421 26776
rect 56227 26816 56285 26817
rect 56227 26776 56236 26816
rect 56276 26776 56285 26816
rect 56227 26775 56285 26776
rect 58827 26816 58869 26825
rect 58827 26776 58828 26816
rect 58868 26776 58869 26816
rect 58827 26767 58869 26776
rect 59019 26816 59061 26825
rect 59019 26776 59020 26816
rect 59060 26776 59061 26816
rect 59019 26767 59061 26776
rect 59107 26816 59165 26817
rect 59107 26776 59116 26816
rect 59156 26776 59165 26816
rect 59107 26775 59165 26776
rect 59491 26816 59549 26817
rect 59491 26776 59500 26816
rect 59540 26776 59549 26816
rect 59491 26775 59549 26776
rect 59787 26816 59829 26825
rect 59787 26776 59788 26816
rect 59828 26776 59829 26816
rect 59787 26767 59829 26776
rect 59883 26816 59925 26825
rect 59883 26776 59884 26816
rect 59924 26776 59925 26816
rect 59883 26767 59925 26776
rect 60739 26816 60797 26817
rect 60739 26776 60748 26816
rect 60788 26776 60797 26816
rect 60739 26775 60797 26776
rect 60939 26816 60981 26825
rect 60939 26776 60940 26816
rect 60980 26776 60981 26816
rect 60939 26767 60981 26776
rect 63819 26816 63861 26825
rect 63819 26776 63820 26816
rect 63860 26776 63861 26816
rect 63819 26767 63861 26776
rect 64011 26816 64053 26825
rect 64011 26776 64012 26816
rect 64052 26776 64053 26816
rect 64011 26767 64053 26776
rect 64099 26816 64157 26817
rect 64099 26776 64108 26816
rect 64148 26776 64157 26816
rect 64099 26775 64157 26776
rect 66787 26816 66845 26817
rect 66787 26776 66796 26816
rect 66836 26776 66845 26816
rect 66787 26775 66845 26776
rect 67651 26816 67709 26817
rect 67651 26776 67660 26816
rect 67700 26776 67709 26816
rect 67651 26775 67709 26776
rect 68331 26816 68373 26825
rect 68331 26776 68332 26816
rect 68372 26776 68373 26816
rect 68331 26767 68373 26776
rect 68523 26816 68565 26825
rect 68523 26776 68524 26816
rect 68564 26776 68565 26816
rect 68523 26767 68565 26776
rect 68611 26816 68669 26817
rect 68611 26776 68620 26816
rect 68660 26776 68669 26816
rect 68611 26775 68669 26776
rect 69195 26816 69237 26825
rect 69195 26776 69196 26816
rect 69236 26776 69237 26816
rect 69195 26767 69237 26776
rect 69571 26816 69629 26817
rect 69571 26776 69580 26816
rect 69620 26776 69629 26816
rect 69571 26775 69629 26776
rect 70435 26816 70493 26817
rect 70435 26776 70444 26816
rect 70484 26776 70493 26816
rect 70435 26775 70493 26776
rect 73035 26816 73077 26825
rect 73035 26776 73036 26816
rect 73076 26776 73077 26816
rect 73411 26812 73420 26852
rect 73460 26812 73469 26852
rect 75435 26851 75477 26860
rect 73411 26811 73469 26812
rect 74275 26816 74333 26817
rect 73035 26767 73077 26776
rect 74275 26776 74284 26816
rect 74324 26776 74333 26816
rect 74275 26775 74333 26776
rect 75627 26816 75669 26825
rect 75627 26776 75628 26816
rect 75668 26776 75669 26816
rect 75627 26767 75669 26776
rect 75723 26816 75765 26825
rect 75723 26776 75724 26816
rect 75764 26776 75765 26816
rect 75723 26767 75765 26776
rect 75819 26816 75861 26825
rect 75819 26776 75820 26816
rect 75860 26776 75861 26816
rect 75819 26767 75861 26776
rect 75915 26816 75957 26825
rect 75915 26776 75916 26816
rect 75956 26776 75957 26816
rect 75915 26767 75957 26776
rect 76195 26816 76253 26817
rect 76195 26776 76204 26816
rect 76244 26776 76253 26816
rect 76195 26775 76253 26776
rect 76491 26816 76533 26825
rect 76491 26776 76492 26816
rect 76532 26776 76533 26816
rect 76491 26767 76533 26776
rect 76587 26816 76629 26825
rect 76587 26776 76588 26816
rect 76628 26776 76629 26816
rect 76587 26767 76629 26776
rect 77443 26816 77501 26817
rect 77443 26776 77452 26816
rect 77492 26776 77501 26816
rect 77443 26775 77501 26776
rect 78307 26816 78365 26817
rect 78307 26776 78316 26816
rect 78356 26776 78365 26816
rect 78307 26775 78365 26776
rect 35691 26732 35733 26741
rect 35691 26692 35692 26732
rect 35732 26692 35733 26732
rect 35691 26683 35733 26692
rect 41451 26732 41493 26741
rect 41451 26692 41452 26732
rect 41492 26692 41493 26732
rect 41451 26683 41493 26692
rect 41739 26732 41781 26741
rect 41739 26692 41740 26732
rect 41780 26692 41781 26732
rect 41739 26683 41781 26692
rect 56619 26732 56661 26741
rect 56619 26692 56620 26732
rect 56660 26692 56661 26732
rect 56619 26683 56661 26692
rect 68043 26732 68085 26741
rect 68043 26692 68044 26732
rect 68084 26692 68085 26732
rect 68043 26683 68085 26692
rect 77067 26732 77109 26741
rect 77067 26692 77068 26732
rect 77108 26692 77109 26732
rect 77067 26683 77109 26692
rect 38083 26648 38141 26649
rect 38083 26608 38092 26648
rect 38132 26608 38141 26648
rect 38083 26607 38141 26608
rect 39723 26648 39765 26657
rect 39723 26608 39724 26648
rect 39764 26608 39765 26648
rect 39723 26599 39765 26608
rect 44131 26648 44189 26649
rect 44131 26608 44140 26648
rect 44180 26608 44189 26648
rect 44131 26607 44189 26608
rect 49507 26648 49565 26649
rect 49507 26608 49516 26648
rect 49556 26608 49565 26648
rect 49507 26607 49565 26608
rect 50187 26648 50229 26657
rect 50187 26608 50188 26648
rect 50228 26608 50229 26648
rect 50187 26599 50229 26608
rect 50659 26648 50717 26649
rect 50659 26608 50668 26648
rect 50708 26608 50717 26648
rect 50659 26607 50717 26608
rect 58539 26648 58581 26657
rect 58539 26608 58540 26648
rect 58580 26608 58581 26648
rect 58539 26599 58581 26608
rect 58915 26648 58973 26649
rect 58915 26608 58924 26648
rect 58964 26608 58973 26648
rect 58915 26607 58973 26608
rect 60555 26648 60597 26657
rect 60555 26608 60556 26648
rect 60596 26608 60597 26648
rect 60555 26599 60597 26608
rect 65635 26648 65693 26649
rect 65635 26608 65644 26648
rect 65684 26608 65693 26648
rect 65635 26607 65693 26608
rect 68419 26648 68477 26649
rect 68419 26608 68428 26648
rect 68468 26608 68477 26648
rect 68419 26607 68477 26608
rect 71587 26648 71645 26649
rect 71587 26608 71596 26648
rect 71636 26608 71645 26648
rect 71587 26607 71645 26608
rect 71979 26648 72021 26657
rect 71979 26608 71980 26648
rect 72020 26608 72021 26648
rect 71979 26599 72021 26608
rect 72171 26648 72213 26657
rect 72171 26608 72172 26648
rect 72212 26608 72213 26648
rect 72171 26599 72213 26608
rect 79459 26648 79517 26649
rect 79459 26608 79468 26648
rect 79508 26608 79517 26648
rect 79459 26607 79517 26608
rect 576 26480 79584 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 76352 26480
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76720 26440 79584 26480
rect 576 26416 79584 26440
rect 35683 26312 35741 26313
rect 35683 26272 35692 26312
rect 35732 26272 35741 26312
rect 35683 26271 35741 26272
rect 39051 26312 39093 26321
rect 39051 26272 39052 26312
rect 39092 26272 39093 26312
rect 39051 26263 39093 26272
rect 40587 26312 40629 26321
rect 40587 26272 40588 26312
rect 40628 26272 40629 26312
rect 40587 26263 40629 26272
rect 40779 26312 40821 26321
rect 40779 26272 40780 26312
rect 40820 26272 40821 26312
rect 40779 26263 40821 26272
rect 41539 26312 41597 26313
rect 41539 26272 41548 26312
rect 41588 26272 41597 26312
rect 41539 26271 41597 26272
rect 46531 26312 46589 26313
rect 46531 26272 46540 26312
rect 46580 26272 46589 26312
rect 46531 26271 46589 26272
rect 52107 26312 52149 26321
rect 52107 26272 52108 26312
rect 52148 26272 52149 26312
rect 52107 26263 52149 26272
rect 56419 26312 56477 26313
rect 56419 26272 56428 26312
rect 56468 26272 56477 26312
rect 56419 26271 56477 26272
rect 59019 26312 59061 26321
rect 59019 26272 59020 26312
rect 59060 26272 59061 26312
rect 59019 26263 59061 26272
rect 61131 26312 61173 26321
rect 61131 26272 61132 26312
rect 61172 26272 61173 26312
rect 61131 26263 61173 26272
rect 67747 26312 67805 26313
rect 67747 26272 67756 26312
rect 67796 26272 67805 26312
rect 67747 26271 67805 26272
rect 69571 26312 69629 26313
rect 69571 26272 69580 26312
rect 69620 26272 69629 26312
rect 69571 26271 69629 26272
rect 70635 26312 70677 26321
rect 70635 26272 70636 26312
rect 70676 26272 70677 26312
rect 70635 26263 70677 26272
rect 74659 26312 74717 26313
rect 74659 26272 74668 26312
rect 74708 26272 74717 26312
rect 74659 26271 74717 26272
rect 76867 26312 76925 26313
rect 76867 26272 76876 26312
rect 76916 26272 76925 26312
rect 76867 26271 76925 26272
rect 35019 26228 35061 26237
rect 35019 26188 35020 26228
rect 35060 26188 35061 26228
rect 35019 26179 35061 26188
rect 48843 26228 48885 26237
rect 48843 26188 48844 26228
rect 48884 26188 48885 26228
rect 48843 26179 48885 26188
rect 51531 26228 51573 26237
rect 51531 26188 51532 26228
rect 51572 26188 51573 26228
rect 51531 26179 51573 26188
rect 55659 26228 55701 26237
rect 55659 26188 55660 26228
rect 55700 26188 55701 26228
rect 55659 26179 55701 26188
rect 61611 26228 61653 26237
rect 61611 26188 61612 26228
rect 61652 26188 61653 26228
rect 61611 26179 61653 26188
rect 64779 26228 64821 26237
rect 64779 26188 64780 26228
rect 64820 26188 64821 26228
rect 64779 26179 64821 26188
rect 71307 26228 71349 26237
rect 71307 26188 71308 26228
rect 71348 26188 71349 26228
rect 71307 26179 71349 26188
rect 71883 26228 71925 26237
rect 71883 26188 71884 26228
rect 71924 26188 71925 26228
rect 71883 26179 71925 26188
rect 75243 26228 75285 26237
rect 75243 26188 75244 26228
rect 75284 26188 75285 26228
rect 75243 26179 75285 26188
rect 33147 26144 33189 26153
rect 33147 26104 33148 26144
rect 33188 26104 33189 26144
rect 33147 26095 33189 26104
rect 33955 26144 34013 26145
rect 33955 26104 33964 26144
rect 34004 26104 34013 26144
rect 33955 26103 34013 26104
rect 34347 26144 34389 26153
rect 34347 26104 34348 26144
rect 34388 26104 34389 26144
rect 34347 26095 34389 26104
rect 34627 26144 34685 26145
rect 34627 26104 34636 26144
rect 34676 26104 34685 26144
rect 34627 26103 34685 26104
rect 34923 26144 34965 26153
rect 34923 26104 34924 26144
rect 34964 26104 34965 26144
rect 34923 26095 34965 26104
rect 35491 26144 35549 26145
rect 35491 26104 35500 26144
rect 35540 26104 35549 26144
rect 35491 26103 35549 26104
rect 35595 26144 35637 26153
rect 35595 26104 35596 26144
rect 35636 26104 35637 26144
rect 35595 26095 35637 26104
rect 35787 26144 35829 26153
rect 35787 26104 35788 26144
rect 35828 26104 35829 26144
rect 35787 26095 35829 26104
rect 39243 26144 39285 26153
rect 39243 26104 39244 26144
rect 39284 26104 39285 26144
rect 39243 26095 39285 26104
rect 39435 26144 39477 26153
rect 39435 26104 39436 26144
rect 39476 26104 39477 26144
rect 39435 26095 39477 26104
rect 39523 26144 39581 26145
rect 39523 26104 39532 26144
rect 39572 26104 39581 26144
rect 39523 26103 39581 26104
rect 39723 26144 39765 26153
rect 39723 26104 39724 26144
rect 39764 26104 39765 26144
rect 39723 26095 39765 26104
rect 39915 26144 39957 26153
rect 39915 26104 39916 26144
rect 39956 26104 39957 26144
rect 39915 26095 39957 26104
rect 40003 26144 40061 26145
rect 40003 26104 40012 26144
rect 40052 26104 40061 26144
rect 40003 26103 40061 26104
rect 41347 26144 41405 26145
rect 41347 26104 41356 26144
rect 41396 26104 41405 26144
rect 41347 26103 41405 26104
rect 41451 26144 41493 26153
rect 41451 26104 41452 26144
rect 41492 26104 41493 26144
rect 41451 26095 41493 26104
rect 41643 26144 41685 26153
rect 41643 26104 41644 26144
rect 41684 26104 41685 26144
rect 41643 26095 41685 26104
rect 43851 26144 43893 26153
rect 43851 26104 43852 26144
rect 43892 26104 43893 26144
rect 43851 26095 43893 26104
rect 44227 26144 44285 26145
rect 44227 26104 44236 26144
rect 44276 26104 44285 26144
rect 44227 26103 44285 26104
rect 45091 26144 45149 26145
rect 45091 26104 45100 26144
rect 45140 26104 45149 26144
rect 45091 26103 45149 26104
rect 46443 26144 46485 26153
rect 46443 26104 46444 26144
rect 46484 26104 46485 26144
rect 46443 26095 46485 26104
rect 46635 26144 46677 26153
rect 46635 26104 46636 26144
rect 46676 26104 46677 26144
rect 46635 26095 46677 26104
rect 46723 26144 46781 26145
rect 46723 26104 46732 26144
rect 46772 26104 46781 26144
rect 46723 26103 46781 26104
rect 47787 26144 47829 26153
rect 47787 26104 47788 26144
rect 47828 26104 47829 26144
rect 47787 26095 47829 26104
rect 48643 26144 48701 26145
rect 48643 26104 48652 26144
rect 48692 26104 48701 26144
rect 48643 26103 48701 26104
rect 49219 26144 49277 26145
rect 49219 26104 49228 26144
rect 49268 26104 49277 26144
rect 49219 26103 49277 26104
rect 50083 26144 50141 26145
rect 50083 26104 50092 26144
rect 50132 26104 50141 26144
rect 50083 26103 50141 26104
rect 51435 26144 51477 26153
rect 51435 26104 51436 26144
rect 51476 26104 51477 26144
rect 51435 26095 51477 26104
rect 51627 26144 51669 26153
rect 51627 26104 51628 26144
rect 51668 26104 51669 26144
rect 51627 26095 51669 26104
rect 51715 26144 51773 26145
rect 51715 26104 51724 26144
rect 51764 26104 51773 26144
rect 51715 26103 51773 26104
rect 52483 26144 52541 26145
rect 52483 26104 52492 26144
rect 52532 26104 52541 26144
rect 52483 26103 52541 26104
rect 52683 26144 52725 26153
rect 52683 26104 52684 26144
rect 52724 26104 52725 26144
rect 52683 26095 52725 26104
rect 54979 26144 55037 26145
rect 54979 26104 54988 26144
rect 55028 26104 55037 26144
rect 54979 26103 55037 26104
rect 55179 26144 55221 26153
rect 55179 26104 55180 26144
rect 55220 26104 55221 26144
rect 55179 26095 55221 26104
rect 55755 26144 55797 26153
rect 55755 26104 55756 26144
rect 55796 26104 55797 26144
rect 55755 26095 55797 26104
rect 56035 26144 56093 26145
rect 56035 26104 56044 26144
rect 56084 26104 56093 26144
rect 56035 26103 56093 26104
rect 56331 26144 56373 26153
rect 56331 26104 56332 26144
rect 56372 26104 56373 26144
rect 56331 26095 56373 26104
rect 56523 26144 56565 26153
rect 56523 26104 56524 26144
rect 56564 26104 56565 26144
rect 56523 26095 56565 26104
rect 56611 26144 56669 26145
rect 56611 26104 56620 26144
rect 56660 26104 56669 26144
rect 56611 26103 56669 26104
rect 56811 26144 56853 26153
rect 56811 26104 56812 26144
rect 56852 26104 56853 26144
rect 56811 26095 56853 26104
rect 57003 26144 57045 26153
rect 57003 26104 57004 26144
rect 57044 26104 57045 26144
rect 57003 26095 57045 26104
rect 57091 26144 57149 26145
rect 57091 26104 57100 26144
rect 57140 26104 57149 26144
rect 57091 26103 57149 26104
rect 58347 26144 58389 26153
rect 58347 26104 58348 26144
rect 58388 26104 58389 26144
rect 58347 26095 58389 26104
rect 58539 26144 58581 26153
rect 58539 26104 58540 26144
rect 58580 26104 58581 26144
rect 58539 26095 58581 26104
rect 58627 26144 58685 26145
rect 58627 26104 58636 26144
rect 58676 26104 58685 26144
rect 59499 26144 59541 26153
rect 58627 26103 58685 26104
rect 59299 26121 59357 26122
rect 59299 26081 59308 26121
rect 59348 26081 59357 26121
rect 59499 26104 59500 26144
rect 59540 26104 59541 26144
rect 59499 26095 59541 26104
rect 59683 26144 59741 26145
rect 59683 26104 59692 26144
rect 59732 26104 59741 26144
rect 59683 26103 59741 26104
rect 59787 26144 59829 26153
rect 59787 26104 59788 26144
rect 59828 26104 59829 26144
rect 59787 26095 59829 26104
rect 59979 26144 60021 26153
rect 59979 26104 59980 26144
rect 60020 26104 60021 26144
rect 59979 26095 60021 26104
rect 61987 26144 62045 26145
rect 61987 26104 61996 26144
rect 62036 26104 62045 26144
rect 61987 26103 62045 26104
rect 62851 26144 62909 26145
rect 62851 26104 62860 26144
rect 62900 26104 62909 26144
rect 62851 26103 62909 26104
rect 64203 26144 64245 26153
rect 64203 26104 64204 26144
rect 64244 26104 64245 26144
rect 64203 26095 64245 26104
rect 64299 26144 64341 26153
rect 64299 26104 64300 26144
rect 64340 26104 64341 26144
rect 64299 26095 64341 26104
rect 64395 26144 64437 26153
rect 64395 26104 64396 26144
rect 64436 26104 64437 26144
rect 64395 26095 64437 26104
rect 64491 26144 64533 26153
rect 64491 26104 64492 26144
rect 64532 26104 64533 26144
rect 64491 26095 64533 26104
rect 64683 26144 64725 26153
rect 64683 26104 64684 26144
rect 64724 26104 64725 26144
rect 64683 26095 64725 26104
rect 64875 26144 64917 26153
rect 64875 26104 64876 26144
rect 64916 26104 64917 26144
rect 64875 26095 64917 26104
rect 64963 26144 65021 26145
rect 64963 26104 64972 26144
rect 65012 26104 65021 26144
rect 64963 26103 65021 26104
rect 65355 26144 65397 26153
rect 65355 26104 65356 26144
rect 65396 26104 65397 26144
rect 65355 26095 65397 26104
rect 65547 26144 65589 26153
rect 65547 26104 65548 26144
rect 65588 26104 65589 26144
rect 65547 26095 65589 26104
rect 65635 26144 65693 26145
rect 65635 26104 65644 26144
rect 65684 26104 65693 26144
rect 65635 26103 65693 26104
rect 67179 26144 67221 26153
rect 67179 26104 67180 26144
rect 67220 26104 67221 26144
rect 67179 26095 67221 26104
rect 67275 26144 67317 26153
rect 67275 26104 67276 26144
rect 67316 26104 67317 26144
rect 67275 26095 67317 26104
rect 67371 26144 67413 26153
rect 67371 26104 67372 26144
rect 67412 26104 67413 26144
rect 67371 26095 67413 26104
rect 67467 26144 67509 26153
rect 67467 26104 67468 26144
rect 67508 26104 67509 26144
rect 67467 26095 67509 26104
rect 67659 26144 67701 26153
rect 67659 26104 67660 26144
rect 67700 26104 67701 26144
rect 67659 26095 67701 26104
rect 67851 26144 67893 26153
rect 67851 26104 67852 26144
rect 67892 26104 67893 26144
rect 67851 26095 67893 26104
rect 67939 26144 67997 26145
rect 67939 26104 67948 26144
rect 67988 26104 67997 26144
rect 67939 26103 67997 26104
rect 68131 26144 68189 26145
rect 68131 26104 68140 26144
rect 68180 26104 68189 26144
rect 68131 26103 68189 26104
rect 68331 26144 68373 26153
rect 68331 26104 68332 26144
rect 68372 26104 68373 26144
rect 68331 26095 68373 26104
rect 69291 26144 69333 26153
rect 69291 26104 69292 26144
rect 69332 26104 69333 26144
rect 69291 26095 69333 26104
rect 69387 26144 69429 26153
rect 69387 26104 69388 26144
rect 69428 26104 69429 26144
rect 69387 26095 69429 26104
rect 69483 26144 69525 26153
rect 69483 26104 69484 26144
rect 69524 26104 69525 26144
rect 69483 26095 69525 26104
rect 70915 26144 70973 26145
rect 70915 26104 70924 26144
rect 70964 26104 70973 26144
rect 70915 26103 70973 26104
rect 71211 26144 71253 26153
rect 71211 26104 71212 26144
rect 71252 26104 71253 26144
rect 71211 26095 71253 26104
rect 71787 26144 71829 26153
rect 71787 26104 71788 26144
rect 71828 26104 71829 26144
rect 71787 26095 71829 26104
rect 71971 26144 72029 26145
rect 71971 26104 71980 26144
rect 72020 26104 72029 26144
rect 71971 26103 72029 26104
rect 74179 26144 74237 26145
rect 74179 26104 74188 26144
rect 74228 26104 74237 26144
rect 74179 26103 74237 26104
rect 74283 26144 74325 26153
rect 74283 26104 74284 26144
rect 74324 26104 74325 26144
rect 74283 26095 74325 26104
rect 74475 26144 74517 26153
rect 74475 26104 74476 26144
rect 74516 26104 74517 26144
rect 74475 26095 74517 26104
rect 74763 26144 74805 26153
rect 74763 26104 74764 26144
rect 74804 26104 74805 26144
rect 74763 26095 74805 26104
rect 74859 26144 74901 26153
rect 74859 26104 74860 26144
rect 74900 26104 74901 26144
rect 74859 26095 74901 26104
rect 74955 26144 74997 26153
rect 74955 26104 74956 26144
rect 74996 26104 74997 26144
rect 74955 26095 74997 26104
rect 75147 26144 75189 26153
rect 75147 26104 75148 26144
rect 75188 26104 75189 26144
rect 75147 26095 75189 26104
rect 75339 26144 75381 26153
rect 75339 26104 75340 26144
rect 75380 26104 75381 26144
rect 75339 26095 75381 26104
rect 75427 26144 75485 26145
rect 75427 26104 75436 26144
rect 75476 26104 75485 26144
rect 75427 26103 75485 26104
rect 76779 26144 76821 26153
rect 76779 26104 76780 26144
rect 76820 26104 76821 26144
rect 76779 26095 76821 26104
rect 76971 26144 77013 26153
rect 76971 26104 76972 26144
rect 77012 26104 77013 26144
rect 76971 26095 77013 26104
rect 77059 26144 77117 26145
rect 77059 26104 77068 26144
rect 77108 26104 77117 26144
rect 77059 26103 77117 26104
rect 59299 26080 59357 26081
rect 643 26060 701 26061
rect 643 26020 652 26060
rect 692 26020 701 26060
rect 643 26019 701 26020
rect 36643 26060 36701 26061
rect 36643 26020 36652 26060
rect 36692 26020 36701 26060
rect 36643 26019 36701 26020
rect 38851 26060 38909 26061
rect 38851 26020 38860 26060
rect 38900 26020 38909 26060
rect 38851 26019 38909 26020
rect 40387 26060 40445 26061
rect 40387 26020 40396 26060
rect 40436 26020 40445 26060
rect 40387 26019 40445 26020
rect 40963 26060 41021 26061
rect 40963 26020 40972 26060
rect 41012 26020 41021 26060
rect 40963 26019 41021 26020
rect 51907 26060 51965 26061
rect 51907 26020 51916 26060
rect 51956 26020 51965 26060
rect 51907 26019 51965 26020
rect 58819 26060 58877 26061
rect 58819 26020 58828 26060
rect 58868 26020 58877 26060
rect 58819 26019 58877 26020
rect 60355 26060 60413 26061
rect 60355 26020 60364 26060
rect 60404 26020 60413 26060
rect 60355 26019 60413 26020
rect 60547 26060 60605 26061
rect 60547 26020 60556 26060
rect 60596 26020 60605 26060
rect 60547 26019 60605 26020
rect 60931 26060 60989 26061
rect 60931 26020 60940 26060
rect 60980 26020 60989 26060
rect 60931 26019 60989 26020
rect 68803 26060 68861 26061
rect 68803 26020 68812 26060
rect 68852 26020 68861 26060
rect 68803 26019 68861 26020
rect 70435 26060 70493 26061
rect 70435 26020 70444 26060
rect 70484 26020 70493 26060
rect 70435 26019 70493 26020
rect 843 25976 885 25985
rect 843 25936 844 25976
rect 884 25936 885 25976
rect 843 25927 885 25936
rect 31939 25976 31997 25977
rect 31939 25936 31948 25976
rect 31988 25936 31997 25976
rect 31939 25935 31997 25936
rect 35299 25976 35357 25977
rect 35299 25936 35308 25976
rect 35348 25936 35357 25976
rect 35299 25935 35357 25936
rect 36267 25976 36309 25985
rect 36267 25936 36268 25976
rect 36308 25936 36309 25976
rect 36267 25927 36309 25936
rect 36843 25976 36885 25985
rect 36843 25936 36844 25976
rect 36884 25936 36885 25976
rect 36843 25927 36885 25936
rect 37707 25976 37749 25985
rect 37707 25936 37708 25976
rect 37748 25936 37749 25976
rect 37707 25927 37749 25936
rect 39723 25976 39765 25985
rect 39723 25936 39724 25976
rect 39764 25936 39765 25976
rect 39723 25927 39765 25936
rect 42219 25976 42261 25985
rect 42219 25936 42220 25976
rect 42260 25936 42261 25976
rect 42219 25927 42261 25936
rect 47403 25976 47445 25985
rect 47403 25936 47404 25976
rect 47444 25936 47445 25976
rect 47403 25927 47445 25936
rect 52875 25976 52917 25985
rect 52875 25936 52876 25976
rect 52916 25936 52917 25976
rect 52875 25927 52917 25936
rect 55083 25976 55125 25985
rect 55083 25936 55084 25976
rect 55124 25936 55125 25976
rect 55083 25927 55125 25936
rect 55363 25976 55421 25977
rect 55363 25936 55372 25976
rect 55412 25936 55421 25976
rect 55363 25935 55421 25936
rect 56811 25976 56853 25985
rect 56811 25936 56812 25976
rect 56852 25936 56853 25976
rect 56811 25927 56853 25936
rect 57963 25976 58005 25985
rect 57963 25936 57964 25976
rect 58004 25936 58005 25976
rect 57963 25927 58005 25936
rect 58347 25976 58389 25985
rect 58347 25936 58348 25976
rect 58388 25936 58389 25976
rect 58347 25927 58389 25936
rect 60171 25976 60213 25985
rect 60171 25936 60172 25976
rect 60212 25936 60213 25976
rect 60171 25927 60213 25936
rect 60747 25976 60789 25985
rect 60747 25936 60748 25976
rect 60788 25936 60789 25976
rect 60747 25927 60789 25936
rect 65355 25976 65397 25985
rect 65355 25936 65356 25976
rect 65396 25936 65397 25976
rect 65355 25927 65397 25936
rect 66411 25976 66453 25985
rect 66411 25936 66412 25976
rect 66452 25936 66453 25976
rect 66411 25927 66453 25936
rect 68619 25976 68661 25985
rect 68619 25936 68620 25976
rect 68660 25936 68661 25976
rect 74475 25976 74517 25985
rect 68619 25927 68661 25936
rect 73419 25934 73461 25943
rect 39243 25892 39285 25901
rect 39243 25852 39244 25892
rect 39284 25852 39285 25892
rect 39243 25843 39285 25852
rect 40587 25892 40629 25901
rect 40587 25852 40588 25892
rect 40628 25852 40629 25892
rect 40587 25843 40629 25852
rect 40779 25892 40821 25901
rect 40779 25852 40780 25892
rect 40820 25852 40821 25892
rect 40779 25843 40821 25852
rect 46243 25892 46301 25893
rect 46243 25852 46252 25892
rect 46292 25852 46301 25892
rect 46243 25851 46301 25852
rect 48363 25892 48405 25901
rect 48363 25852 48364 25892
rect 48404 25852 48405 25892
rect 48363 25843 48405 25852
rect 51235 25892 51293 25893
rect 51235 25852 51244 25892
rect 51284 25852 51293 25892
rect 51235 25851 51293 25852
rect 52107 25892 52149 25901
rect 52107 25852 52108 25892
rect 52148 25852 52149 25892
rect 52107 25843 52149 25852
rect 52587 25892 52629 25901
rect 52587 25852 52588 25892
rect 52628 25852 52629 25892
rect 52587 25843 52629 25852
rect 59019 25892 59061 25901
rect 59019 25852 59020 25892
rect 59060 25852 59061 25892
rect 59019 25843 59061 25852
rect 59403 25892 59445 25901
rect 59403 25852 59404 25892
rect 59444 25852 59445 25892
rect 59403 25843 59445 25852
rect 59979 25892 60021 25901
rect 59979 25852 59980 25892
rect 60020 25852 60021 25892
rect 59979 25843 60021 25852
rect 64003 25892 64061 25893
rect 64003 25852 64012 25892
rect 64052 25852 64061 25892
rect 64003 25851 64061 25852
rect 68235 25892 68277 25901
rect 73419 25894 73420 25934
rect 73460 25894 73461 25934
rect 74475 25936 74476 25976
rect 74516 25936 74517 25976
rect 74475 25927 74517 25936
rect 68235 25852 68236 25892
rect 68276 25852 68277 25892
rect 68235 25843 68277 25852
rect 71587 25892 71645 25893
rect 71587 25852 71596 25892
rect 71636 25852 71645 25892
rect 73419 25885 73461 25894
rect 71587 25851 71645 25852
rect 576 25724 79584 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 75112 25724
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75480 25684 79584 25724
rect 576 25660 79584 25684
rect 34731 25556 34773 25565
rect 34731 25516 34732 25556
rect 34772 25516 34773 25556
rect 34731 25507 34773 25516
rect 35403 25556 35445 25565
rect 35403 25516 35404 25556
rect 35444 25516 35445 25556
rect 35403 25507 35445 25516
rect 35691 25556 35733 25565
rect 35691 25516 35692 25556
rect 35732 25516 35733 25556
rect 35691 25507 35733 25516
rect 40395 25556 40437 25565
rect 40395 25516 40396 25556
rect 40436 25516 40437 25556
rect 40395 25507 40437 25516
rect 40875 25556 40917 25565
rect 40875 25516 40876 25556
rect 40916 25516 40917 25556
rect 40875 25507 40917 25516
rect 44043 25556 44085 25565
rect 44043 25516 44044 25556
rect 44084 25516 44085 25556
rect 44043 25507 44085 25516
rect 54787 25556 54845 25557
rect 54787 25516 54796 25556
rect 54836 25516 54845 25556
rect 54787 25515 54845 25516
rect 67747 25556 67805 25557
rect 67747 25516 67756 25556
rect 67796 25516 67805 25556
rect 67747 25515 67805 25516
rect 75619 25556 75677 25557
rect 75619 25516 75628 25556
rect 75668 25516 75677 25556
rect 75619 25515 75677 25516
rect 30315 25472 30357 25481
rect 30315 25432 30316 25472
rect 30356 25432 30357 25472
rect 30315 25423 30357 25432
rect 32715 25472 32757 25481
rect 32715 25432 32716 25472
rect 32756 25432 32757 25472
rect 32715 25423 32757 25432
rect 41355 25472 41397 25481
rect 41355 25432 41356 25472
rect 41396 25432 41397 25472
rect 41355 25423 41397 25432
rect 42795 25472 42837 25481
rect 42795 25432 42796 25472
rect 42836 25432 42837 25472
rect 42795 25423 42837 25432
rect 43851 25472 43893 25481
rect 43851 25432 43852 25472
rect 43892 25432 43893 25472
rect 43851 25423 43893 25432
rect 46347 25472 46389 25481
rect 46347 25432 46348 25472
rect 46388 25432 46389 25472
rect 46347 25423 46389 25432
rect 51427 25472 51485 25473
rect 51427 25432 51436 25472
rect 51476 25432 51485 25472
rect 51427 25431 51485 25432
rect 55563 25472 55605 25481
rect 55563 25432 55564 25472
rect 55604 25432 55605 25472
rect 55563 25423 55605 25432
rect 63811 25472 63869 25473
rect 63811 25432 63820 25472
rect 63860 25432 63869 25472
rect 63811 25431 63869 25432
rect 73027 25472 73085 25473
rect 73027 25432 73036 25472
rect 73076 25432 73085 25472
rect 73027 25431 73085 25432
rect 75915 25472 75957 25481
rect 75915 25432 75916 25472
rect 75956 25432 75957 25472
rect 75915 25423 75957 25432
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 40675 25388 40733 25389
rect 40675 25348 40684 25388
rect 40724 25348 40733 25388
rect 40675 25347 40733 25348
rect 31947 25304 31989 25313
rect 31947 25264 31948 25304
rect 31988 25264 31989 25304
rect 31947 25255 31989 25264
rect 32043 25304 32085 25313
rect 32043 25264 32044 25304
rect 32084 25264 32085 25304
rect 32043 25255 32085 25264
rect 32139 25304 32181 25313
rect 32139 25264 32140 25304
rect 32180 25264 32181 25304
rect 32139 25255 32181 25264
rect 33195 25304 33237 25313
rect 33195 25264 33196 25304
rect 33236 25264 33237 25304
rect 33195 25255 33237 25264
rect 33387 25304 33429 25313
rect 33387 25264 33388 25304
rect 33428 25264 33429 25304
rect 33387 25255 33429 25264
rect 33475 25304 33533 25305
rect 33475 25264 33484 25304
rect 33524 25264 33533 25304
rect 33475 25263 33533 25264
rect 34251 25304 34293 25313
rect 34251 25264 34252 25304
rect 34292 25264 34293 25304
rect 34251 25255 34293 25264
rect 34347 25304 34389 25313
rect 34347 25264 34348 25304
rect 34388 25264 34389 25304
rect 34347 25255 34389 25264
rect 34443 25304 34485 25313
rect 34443 25264 34444 25304
rect 34484 25264 34485 25304
rect 34443 25255 34485 25264
rect 34539 25304 34581 25313
rect 34539 25264 34540 25304
rect 34580 25264 34581 25304
rect 34539 25255 34581 25264
rect 34731 25304 34773 25313
rect 34731 25264 34732 25304
rect 34772 25264 34773 25304
rect 34731 25255 34773 25264
rect 34923 25304 34965 25313
rect 34923 25264 34924 25304
rect 34964 25264 34965 25304
rect 34923 25255 34965 25264
rect 35011 25304 35069 25305
rect 35011 25264 35020 25304
rect 35060 25264 35069 25304
rect 35011 25263 35069 25264
rect 35307 25304 35349 25313
rect 35307 25264 35308 25304
rect 35348 25264 35349 25304
rect 35307 25255 35349 25264
rect 35491 25304 35549 25305
rect 35491 25264 35500 25304
rect 35540 25264 35549 25304
rect 35491 25263 35549 25264
rect 35691 25304 35733 25313
rect 35691 25264 35692 25304
rect 35732 25264 35733 25304
rect 35691 25255 35733 25264
rect 35883 25304 35925 25313
rect 35883 25264 35884 25304
rect 35924 25264 35925 25304
rect 35883 25255 35925 25264
rect 35971 25304 36029 25305
rect 35971 25264 35980 25304
rect 36020 25264 36029 25304
rect 35971 25263 36029 25264
rect 36355 25304 36413 25305
rect 36355 25264 36364 25304
rect 36404 25264 36413 25304
rect 36355 25263 36413 25264
rect 37227 25304 37269 25313
rect 37227 25264 37228 25304
rect 37268 25264 37269 25304
rect 37227 25255 37269 25264
rect 37603 25304 37661 25305
rect 37603 25264 37612 25304
rect 37652 25264 37661 25304
rect 37603 25263 37661 25264
rect 38467 25304 38525 25305
rect 38467 25264 38476 25304
rect 38516 25264 38525 25304
rect 38467 25263 38525 25264
rect 39819 25304 39861 25313
rect 39819 25264 39820 25304
rect 39860 25264 39861 25304
rect 39819 25255 39861 25264
rect 39915 25304 39957 25313
rect 39915 25264 39916 25304
rect 39956 25264 39957 25304
rect 39915 25255 39957 25264
rect 40011 25304 40053 25313
rect 40011 25264 40012 25304
rect 40052 25264 40053 25304
rect 40011 25255 40053 25264
rect 40107 25304 40149 25313
rect 40107 25264 40108 25304
rect 40148 25264 40149 25304
rect 40107 25255 40149 25264
rect 40299 25304 40341 25313
rect 40299 25264 40300 25304
rect 40340 25264 40341 25304
rect 40299 25255 40341 25264
rect 40483 25304 40541 25305
rect 40483 25264 40492 25304
rect 40532 25264 40541 25304
rect 40483 25263 40541 25264
rect 44043 25304 44085 25313
rect 44043 25264 44044 25304
rect 44084 25264 44085 25304
rect 44043 25255 44085 25264
rect 44235 25304 44277 25313
rect 44235 25264 44236 25304
rect 44276 25264 44277 25304
rect 44235 25255 44277 25264
rect 44323 25304 44381 25305
rect 44323 25264 44332 25304
rect 44372 25264 44381 25304
rect 44323 25263 44381 25264
rect 44619 25304 44661 25313
rect 44619 25264 44620 25304
rect 44660 25264 44661 25304
rect 44619 25255 44661 25264
rect 44715 25304 44757 25313
rect 44715 25264 44716 25304
rect 44756 25264 44757 25304
rect 44715 25255 44757 25264
rect 44811 25304 44853 25313
rect 44811 25264 44812 25304
rect 44852 25264 44853 25304
rect 44811 25255 44853 25264
rect 45955 25304 46013 25305
rect 45955 25264 45964 25304
rect 46004 25264 46013 25304
rect 45955 25263 46013 25264
rect 46251 25304 46293 25313
rect 46251 25264 46252 25304
rect 46292 25264 46293 25304
rect 46251 25255 46293 25264
rect 46435 25304 46493 25305
rect 46435 25264 46444 25304
rect 46484 25264 46493 25304
rect 46435 25263 46493 25264
rect 46731 25304 46773 25313
rect 46731 25264 46732 25304
rect 46772 25264 46773 25304
rect 46731 25255 46773 25264
rect 46915 25304 46973 25305
rect 46915 25264 46924 25304
rect 46964 25264 46973 25304
rect 46915 25263 46973 25264
rect 47491 25304 47549 25305
rect 47491 25264 47500 25304
rect 47540 25264 47549 25304
rect 47491 25263 47549 25264
rect 48355 25304 48413 25305
rect 48355 25264 48364 25304
rect 48404 25264 48413 25304
rect 48355 25263 48413 25264
rect 50571 25304 50613 25313
rect 50571 25264 50572 25304
rect 50612 25264 50613 25304
rect 50571 25255 50613 25264
rect 50667 25304 50709 25313
rect 50667 25264 50668 25304
rect 50708 25264 50709 25304
rect 50667 25255 50709 25264
rect 50763 25304 50805 25313
rect 50763 25264 50764 25304
rect 50804 25264 50805 25304
rect 50763 25255 50805 25264
rect 50859 25304 50901 25313
rect 50859 25264 50860 25304
rect 50900 25264 50901 25304
rect 50859 25255 50901 25264
rect 51043 25304 51101 25305
rect 51043 25264 51052 25304
rect 51092 25264 51101 25304
rect 51043 25263 51101 25264
rect 51243 25304 51285 25313
rect 51243 25264 51244 25304
rect 51284 25264 51285 25304
rect 51243 25255 51285 25264
rect 51723 25304 51765 25313
rect 51723 25264 51724 25304
rect 51764 25264 51765 25304
rect 51723 25255 51765 25264
rect 51819 25304 51861 25313
rect 51819 25264 51820 25304
rect 51860 25264 51861 25304
rect 51819 25255 51861 25264
rect 52099 25304 52157 25305
rect 52099 25264 52108 25304
rect 52148 25264 52157 25304
rect 52099 25263 52157 25264
rect 52771 25304 52829 25305
rect 52771 25264 52780 25304
rect 52820 25264 52829 25304
rect 52771 25263 52829 25264
rect 53635 25304 53693 25305
rect 53635 25264 53644 25304
rect 53684 25264 53693 25304
rect 53635 25263 53693 25264
rect 55747 25304 55805 25305
rect 55747 25264 55756 25304
rect 55796 25264 55805 25304
rect 55747 25263 55805 25264
rect 55947 25304 55989 25313
rect 55947 25264 55948 25304
rect 55988 25264 55989 25304
rect 55947 25255 55989 25264
rect 57483 25304 57525 25313
rect 57483 25264 57484 25304
rect 57524 25264 57525 25304
rect 57483 25255 57525 25264
rect 57859 25304 57917 25305
rect 57859 25264 57868 25304
rect 57908 25264 57917 25304
rect 57859 25263 57917 25264
rect 58723 25304 58781 25305
rect 58723 25264 58732 25304
rect 58772 25264 58781 25304
rect 58723 25263 58781 25264
rect 60171 25304 60213 25313
rect 60171 25264 60172 25304
rect 60212 25264 60213 25304
rect 60171 25255 60213 25264
rect 60547 25304 60605 25305
rect 60547 25264 60556 25304
rect 60596 25264 60605 25304
rect 60547 25263 60605 25264
rect 61411 25304 61469 25305
rect 61411 25264 61420 25304
rect 61460 25264 61469 25304
rect 61411 25263 61469 25264
rect 63139 25304 63197 25305
rect 63139 25264 63148 25304
rect 63188 25264 63197 25304
rect 63139 25263 63197 25264
rect 63435 25304 63477 25313
rect 63435 25264 63436 25304
rect 63476 25264 63477 25304
rect 63435 25255 63477 25264
rect 63531 25304 63573 25313
rect 63531 25264 63532 25304
rect 63572 25264 63573 25304
rect 63531 25255 63573 25264
rect 64387 25304 64445 25305
rect 64387 25264 64396 25304
rect 64436 25264 64445 25304
rect 64387 25263 64445 25264
rect 65251 25304 65309 25305
rect 65251 25264 65260 25304
rect 65300 25264 65309 25304
rect 65251 25263 65309 25264
rect 67075 25304 67133 25305
rect 67075 25264 67084 25304
rect 67124 25264 67133 25304
rect 67075 25263 67133 25264
rect 67371 25304 67413 25313
rect 67371 25264 67372 25304
rect 67412 25264 67413 25304
rect 67371 25255 67413 25264
rect 67467 25304 67509 25313
rect 67467 25264 67468 25304
rect 67508 25264 67509 25304
rect 69187 25304 69245 25305
rect 67467 25255 67509 25264
rect 68323 25291 68381 25292
rect 68323 25251 68332 25291
rect 68372 25251 68381 25291
rect 69187 25264 69196 25304
rect 69236 25264 69245 25304
rect 69187 25263 69245 25264
rect 71011 25304 71069 25305
rect 71011 25264 71020 25304
rect 71060 25264 71069 25304
rect 71011 25263 71069 25264
rect 71875 25304 71933 25305
rect 71875 25264 71884 25304
rect 71924 25264 71933 25304
rect 71875 25263 71933 25264
rect 73227 25304 73269 25313
rect 73227 25264 73228 25304
rect 73268 25264 73269 25304
rect 73227 25255 73269 25264
rect 73603 25304 73661 25305
rect 73603 25264 73612 25304
rect 73652 25264 73661 25304
rect 73603 25263 73661 25264
rect 74467 25304 74525 25305
rect 74467 25264 74476 25304
rect 74516 25264 74525 25304
rect 74467 25263 74525 25264
rect 75811 25304 75869 25305
rect 75811 25264 75820 25304
rect 75860 25264 75869 25304
rect 75811 25263 75869 25264
rect 76011 25304 76053 25313
rect 76011 25264 76012 25304
rect 76052 25264 76053 25304
rect 76011 25255 76053 25264
rect 76203 25304 76245 25313
rect 76203 25264 76204 25304
rect 76244 25264 76245 25304
rect 76203 25255 76245 25264
rect 76395 25304 76437 25313
rect 76395 25264 76396 25304
rect 76436 25264 76437 25304
rect 76395 25255 76437 25264
rect 76483 25304 76541 25305
rect 76483 25264 76492 25304
rect 76532 25264 76541 25304
rect 76483 25263 76541 25264
rect 77059 25304 77117 25305
rect 77059 25264 77068 25304
rect 77108 25264 77117 25304
rect 77059 25263 77117 25264
rect 77923 25304 77981 25305
rect 77923 25264 77932 25304
rect 77972 25264 77981 25304
rect 77923 25263 77981 25264
rect 68323 25250 68381 25251
rect 46827 25220 46869 25229
rect 46827 25180 46828 25220
rect 46868 25180 46869 25220
rect 46827 25171 46869 25180
rect 47115 25220 47157 25229
rect 47115 25180 47116 25220
rect 47156 25180 47157 25220
rect 47115 25171 47157 25180
rect 51147 25220 51189 25229
rect 51147 25180 51148 25220
rect 51188 25180 51189 25220
rect 51147 25171 51189 25180
rect 52395 25220 52437 25229
rect 52395 25180 52396 25220
rect 52436 25180 52437 25220
rect 52395 25171 52437 25180
rect 55851 25220 55893 25229
rect 55851 25180 55852 25220
rect 55892 25180 55893 25220
rect 55851 25171 55893 25180
rect 64011 25220 64053 25229
rect 64011 25180 64012 25220
rect 64052 25180 64053 25220
rect 64011 25171 64053 25180
rect 67947 25220 67989 25229
rect 67947 25180 67948 25220
rect 67988 25180 67989 25220
rect 67947 25171 67989 25180
rect 70635 25220 70677 25229
rect 70635 25180 70636 25220
rect 70676 25180 70677 25220
rect 70635 25171 70677 25180
rect 76299 25220 76341 25229
rect 76299 25180 76300 25220
rect 76340 25180 76341 25220
rect 76299 25171 76341 25180
rect 76683 25220 76725 25229
rect 76683 25180 76684 25220
rect 76724 25180 76725 25220
rect 76683 25171 76725 25180
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 32227 25136 32285 25137
rect 32227 25096 32236 25136
rect 32276 25096 32285 25136
rect 32227 25095 32285 25096
rect 33283 25136 33341 25137
rect 33283 25096 33292 25136
rect 33332 25096 33341 25136
rect 33283 25095 33341 25096
rect 39619 25136 39677 25137
rect 39619 25096 39628 25136
rect 39668 25096 39677 25136
rect 39619 25095 39677 25096
rect 40875 25136 40917 25145
rect 40875 25096 40876 25136
rect 40916 25096 40917 25136
rect 40875 25087 40917 25096
rect 44515 25136 44573 25137
rect 44515 25096 44524 25136
rect 44564 25096 44573 25136
rect 44515 25095 44573 25096
rect 49507 25136 49565 25137
rect 49507 25096 49516 25136
rect 49556 25096 49565 25136
rect 49507 25095 49565 25096
rect 54787 25136 54845 25137
rect 54787 25096 54796 25136
rect 54836 25096 54845 25136
rect 54787 25095 54845 25096
rect 59875 25136 59933 25137
rect 59875 25096 59884 25136
rect 59924 25096 59933 25136
rect 59875 25095 59933 25096
rect 62563 25136 62621 25137
rect 62563 25096 62572 25136
rect 62612 25096 62621 25136
rect 62563 25095 62621 25096
rect 66403 25136 66461 25137
rect 66403 25096 66412 25136
rect 66452 25096 66461 25136
rect 66403 25095 66461 25096
rect 70339 25136 70397 25137
rect 70339 25096 70348 25136
rect 70388 25096 70397 25136
rect 70339 25095 70397 25096
rect 75619 25136 75677 25137
rect 75619 25096 75628 25136
rect 75668 25096 75677 25136
rect 75619 25095 75677 25096
rect 79075 25136 79133 25137
rect 79075 25096 79084 25136
rect 79124 25096 79133 25136
rect 79075 25095 79133 25096
rect 576 24968 79584 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 76352 24968
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76720 24928 79584 24968
rect 576 24904 79584 24928
rect 37507 24800 37565 24801
rect 37507 24760 37516 24800
rect 37556 24760 37565 24800
rect 37507 24759 37565 24760
rect 44995 24800 45053 24801
rect 44995 24760 45004 24800
rect 45044 24760 45053 24800
rect 44995 24759 45053 24760
rect 50187 24800 50229 24809
rect 50187 24760 50188 24800
rect 50228 24760 50229 24800
rect 50187 24751 50229 24760
rect 58339 24800 58397 24801
rect 58339 24760 58348 24800
rect 58388 24760 58397 24800
rect 58339 24759 58397 24760
rect 58923 24800 58965 24809
rect 58923 24760 58924 24800
rect 58964 24760 58965 24800
rect 58923 24751 58965 24760
rect 60459 24800 60501 24809
rect 60459 24760 60460 24800
rect 60500 24760 60501 24800
rect 60459 24751 60501 24760
rect 64003 24800 64061 24801
rect 64003 24760 64012 24800
rect 64052 24760 64061 24800
rect 64003 24759 64061 24760
rect 67747 24800 67805 24801
rect 67747 24760 67756 24800
rect 67796 24760 67805 24800
rect 67747 24759 67805 24760
rect 70819 24800 70877 24801
rect 70819 24760 70828 24800
rect 70868 24760 70877 24800
rect 70819 24759 70877 24760
rect 74371 24800 74429 24801
rect 74371 24760 74380 24800
rect 74420 24760 74429 24800
rect 74371 24759 74429 24760
rect 29835 24716 29877 24725
rect 29835 24676 29836 24716
rect 29876 24676 29877 24716
rect 29835 24667 29877 24676
rect 32523 24716 32565 24725
rect 32523 24676 32524 24716
rect 32564 24676 32565 24716
rect 32523 24667 32565 24676
rect 46443 24716 46485 24725
rect 46443 24676 46444 24716
rect 46484 24676 46485 24716
rect 59403 24716 59445 24725
rect 46443 24667 46485 24676
rect 50379 24674 50421 24683
rect 30211 24632 30269 24633
rect 30211 24592 30220 24632
rect 30260 24592 30269 24632
rect 30211 24591 30269 24592
rect 31075 24632 31133 24633
rect 31075 24592 31084 24632
rect 31124 24592 31133 24632
rect 31075 24591 31133 24592
rect 32427 24632 32469 24641
rect 32427 24592 32428 24632
rect 32468 24592 32469 24632
rect 32427 24583 32469 24592
rect 32619 24632 32661 24641
rect 32619 24592 32620 24632
rect 32660 24592 32661 24632
rect 32619 24583 32661 24592
rect 32707 24632 32765 24633
rect 32707 24592 32716 24632
rect 32756 24592 32765 24632
rect 32707 24591 32765 24592
rect 35115 24632 35157 24641
rect 35115 24592 35116 24632
rect 35156 24592 35157 24632
rect 35115 24583 35157 24592
rect 35491 24632 35549 24633
rect 35491 24592 35500 24632
rect 35540 24592 35549 24632
rect 35491 24591 35549 24592
rect 36355 24632 36413 24633
rect 36355 24592 36364 24632
rect 36404 24592 36413 24632
rect 36355 24591 36413 24592
rect 39523 24632 39581 24633
rect 39523 24592 39532 24632
rect 39572 24592 39581 24632
rect 39523 24591 39581 24592
rect 39819 24632 39861 24641
rect 39819 24592 39820 24632
rect 39860 24592 39861 24632
rect 39819 24583 39861 24592
rect 39915 24632 39957 24641
rect 39915 24592 39916 24632
rect 39956 24592 39957 24632
rect 39915 24583 39957 24592
rect 40395 24632 40437 24641
rect 40395 24592 40396 24632
rect 40436 24592 40437 24632
rect 40395 24583 40437 24592
rect 40587 24632 40629 24641
rect 40587 24592 40588 24632
rect 40628 24592 40629 24632
rect 40587 24583 40629 24592
rect 40675 24632 40733 24633
rect 40675 24592 40684 24632
rect 40724 24592 40733 24632
rect 40675 24591 40733 24592
rect 40867 24632 40925 24633
rect 40867 24592 40876 24632
rect 40916 24592 40925 24632
rect 40867 24591 40925 24592
rect 40971 24632 41013 24641
rect 40971 24592 40972 24632
rect 41012 24592 41013 24632
rect 40971 24583 41013 24592
rect 41067 24632 41109 24641
rect 41067 24592 41068 24632
rect 41108 24592 41109 24632
rect 41067 24583 41109 24592
rect 42315 24632 42357 24641
rect 42315 24592 42316 24632
rect 42356 24592 42357 24632
rect 42315 24583 42357 24592
rect 42691 24632 42749 24633
rect 42691 24592 42700 24632
rect 42740 24592 42749 24632
rect 42691 24591 42749 24592
rect 43555 24632 43613 24633
rect 43555 24592 43564 24632
rect 43604 24592 43613 24632
rect 43555 24591 43613 24592
rect 44907 24632 44949 24641
rect 44907 24592 44908 24632
rect 44948 24592 44949 24632
rect 44907 24583 44949 24592
rect 45099 24632 45141 24641
rect 45099 24592 45100 24632
rect 45140 24592 45141 24632
rect 45099 24583 45141 24592
rect 45187 24632 45245 24633
rect 45187 24592 45196 24632
rect 45236 24592 45245 24632
rect 45187 24591 45245 24592
rect 46539 24632 46581 24641
rect 46539 24592 46540 24632
rect 46580 24592 46581 24632
rect 46539 24583 46581 24592
rect 46819 24632 46877 24633
rect 46819 24592 46828 24632
rect 46868 24592 46877 24632
rect 46819 24591 46877 24592
rect 47115 24632 47157 24641
rect 47115 24592 47116 24632
rect 47156 24592 47157 24632
rect 47115 24583 47157 24592
rect 47307 24632 47349 24641
rect 50379 24634 50380 24674
rect 50420 24634 50421 24674
rect 59403 24676 59404 24716
rect 59444 24676 59445 24716
rect 59403 24667 59445 24676
rect 60171 24716 60213 24725
rect 60171 24676 60172 24716
rect 60212 24676 60213 24716
rect 60171 24667 60213 24676
rect 64491 24716 64533 24725
rect 64491 24676 64492 24716
rect 64532 24676 64533 24716
rect 64491 24667 64533 24676
rect 68235 24716 68277 24725
rect 68235 24676 68236 24716
rect 68276 24676 68277 24716
rect 68235 24667 68277 24676
rect 75819 24716 75861 24725
rect 75819 24676 75820 24716
rect 75860 24676 75861 24716
rect 75819 24667 75861 24676
rect 76587 24716 76629 24725
rect 76587 24676 76588 24716
rect 76628 24676 76629 24716
rect 76587 24667 76629 24676
rect 47307 24592 47308 24632
rect 47348 24592 47349 24632
rect 47307 24583 47349 24592
rect 47395 24632 47453 24633
rect 47395 24592 47404 24632
rect 47444 24592 47453 24632
rect 50379 24625 50421 24634
rect 50571 24632 50613 24641
rect 47395 24591 47453 24592
rect 50571 24592 50572 24632
rect 50612 24592 50613 24632
rect 50571 24583 50613 24592
rect 50659 24632 50717 24633
rect 50659 24592 50668 24632
rect 50708 24592 50717 24632
rect 50659 24591 50717 24592
rect 52107 24632 52149 24641
rect 52107 24592 52108 24632
rect 52148 24592 52149 24632
rect 52107 24583 52149 24592
rect 52299 24632 52341 24641
rect 52299 24592 52300 24632
rect 52340 24592 52341 24632
rect 52299 24583 52341 24592
rect 52387 24632 52445 24633
rect 52387 24592 52396 24632
rect 52436 24592 52445 24632
rect 52387 24591 52445 24592
rect 55083 24632 55125 24641
rect 55083 24592 55084 24632
rect 55124 24592 55125 24632
rect 55083 24583 55125 24592
rect 55459 24632 55517 24633
rect 55459 24592 55468 24632
rect 55508 24592 55517 24632
rect 55459 24591 55517 24592
rect 56323 24632 56381 24633
rect 56323 24592 56332 24632
rect 56372 24592 56381 24632
rect 56323 24591 56381 24592
rect 58059 24632 58101 24641
rect 58059 24592 58060 24632
rect 58100 24592 58101 24632
rect 58059 24583 58101 24592
rect 58155 24632 58197 24641
rect 58155 24592 58156 24632
rect 58196 24592 58197 24632
rect 58155 24583 58197 24592
rect 58251 24632 58293 24641
rect 58251 24592 58252 24632
rect 58292 24592 58293 24632
rect 58251 24583 58293 24592
rect 59499 24632 59541 24641
rect 59499 24592 59500 24632
rect 59540 24592 59541 24632
rect 59499 24583 59541 24592
rect 59779 24632 59837 24633
rect 59779 24592 59788 24632
rect 59828 24592 59837 24632
rect 59779 24591 59837 24592
rect 60075 24632 60117 24641
rect 60075 24592 60076 24632
rect 60116 24592 60117 24632
rect 60075 24583 60117 24592
rect 60259 24632 60317 24633
rect 60259 24592 60268 24632
rect 60308 24592 60317 24632
rect 60259 24591 60317 24592
rect 63523 24632 63581 24633
rect 63523 24592 63532 24632
rect 63572 24592 63581 24632
rect 63523 24591 63581 24592
rect 63627 24632 63669 24641
rect 63627 24592 63628 24632
rect 63668 24592 63669 24632
rect 63627 24583 63669 24592
rect 63723 24632 63765 24641
rect 63723 24592 63724 24632
rect 63764 24592 63765 24632
rect 63723 24583 63765 24592
rect 63915 24632 63957 24641
rect 63915 24592 63916 24632
rect 63956 24592 63957 24632
rect 63915 24583 63957 24592
rect 64107 24632 64149 24641
rect 64107 24592 64108 24632
rect 64148 24592 64149 24632
rect 64107 24583 64149 24592
rect 64195 24632 64253 24633
rect 64195 24592 64204 24632
rect 64244 24592 64253 24632
rect 64195 24591 64253 24592
rect 64387 24632 64445 24633
rect 64387 24592 64396 24632
rect 64436 24592 64445 24632
rect 64387 24591 64445 24592
rect 64587 24632 64629 24641
rect 64587 24592 64588 24632
rect 64628 24592 64629 24632
rect 64587 24583 64629 24592
rect 67659 24632 67701 24641
rect 67659 24592 67660 24632
rect 67700 24592 67701 24632
rect 67659 24583 67701 24592
rect 67851 24632 67893 24641
rect 67851 24592 67852 24632
rect 67892 24592 67893 24632
rect 67851 24583 67893 24592
rect 67939 24632 67997 24633
rect 67939 24592 67948 24632
rect 67988 24592 67997 24632
rect 67939 24591 67997 24592
rect 68131 24632 68189 24633
rect 68131 24592 68140 24632
rect 68180 24592 68189 24632
rect 68131 24591 68189 24592
rect 68331 24632 68373 24641
rect 68331 24592 68332 24632
rect 68372 24592 68373 24632
rect 68331 24583 68373 24592
rect 70731 24632 70773 24641
rect 70731 24592 70732 24632
rect 70772 24592 70773 24632
rect 70731 24583 70773 24592
rect 70923 24632 70965 24641
rect 70923 24592 70924 24632
rect 70964 24592 70965 24632
rect 70923 24583 70965 24592
rect 71011 24632 71069 24633
rect 71011 24592 71020 24632
rect 71060 24592 71069 24632
rect 71011 24591 71069 24592
rect 71587 24632 71645 24633
rect 71587 24592 71596 24632
rect 71636 24592 71645 24632
rect 71587 24591 71645 24592
rect 71691 24632 71733 24641
rect 71691 24592 71692 24632
rect 71732 24592 71733 24632
rect 71691 24583 71733 24592
rect 71787 24632 71829 24641
rect 71787 24592 71788 24632
rect 71828 24592 71829 24632
rect 71787 24583 71829 24592
rect 74283 24632 74325 24641
rect 74283 24592 74284 24632
rect 74324 24592 74325 24632
rect 74283 24583 74325 24592
rect 74475 24632 74517 24641
rect 74475 24592 74476 24632
rect 74516 24592 74517 24632
rect 74475 24583 74517 24592
rect 74563 24632 74621 24633
rect 74563 24592 74572 24632
rect 74612 24592 74621 24632
rect 74563 24591 74621 24592
rect 75427 24632 75485 24633
rect 75427 24592 75436 24632
rect 75476 24592 75485 24632
rect 75427 24591 75485 24592
rect 75723 24632 75765 24641
rect 75723 24592 75724 24632
rect 75764 24592 75765 24632
rect 75723 24583 75765 24592
rect 76483 24632 76541 24633
rect 76483 24592 76492 24632
rect 76532 24592 76541 24632
rect 76483 24591 76541 24592
rect 76683 24632 76725 24641
rect 76683 24592 76684 24632
rect 76724 24592 76725 24632
rect 76683 24583 76725 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 39043 24548 39101 24549
rect 39043 24508 39052 24548
rect 39092 24508 39101 24548
rect 39043 24507 39101 24508
rect 49987 24548 50045 24549
rect 49987 24508 49996 24548
rect 50036 24508 50045 24548
rect 49987 24507 50045 24508
rect 51331 24548 51389 24549
rect 51331 24508 51340 24548
rect 51380 24508 51389 24548
rect 51331 24507 51389 24508
rect 57483 24548 57525 24557
rect 57483 24508 57484 24548
rect 57524 24508 57525 24548
rect 57483 24499 57525 24508
rect 58723 24548 58781 24549
rect 58723 24508 58732 24548
rect 58772 24508 58781 24548
rect 58723 24507 58781 24508
rect 60643 24548 60701 24549
rect 60643 24508 60652 24548
rect 60692 24508 60701 24548
rect 60643 24507 60701 24508
rect 40195 24464 40253 24465
rect 40195 24424 40204 24464
rect 40244 24424 40253 24464
rect 40195 24423 40253 24424
rect 46147 24464 46205 24465
rect 46147 24424 46156 24464
rect 46196 24424 46205 24464
rect 46147 24423 46205 24424
rect 47115 24464 47157 24473
rect 47115 24424 47116 24464
rect 47156 24424 47157 24464
rect 47115 24415 47157 24424
rect 47595 24464 47637 24473
rect 47595 24424 47596 24464
rect 47636 24424 47637 24464
rect 47595 24415 47637 24424
rect 48459 24464 48501 24473
rect 48459 24424 48460 24464
rect 48500 24424 48501 24464
rect 48459 24415 48501 24424
rect 51147 24464 51189 24473
rect 51147 24424 51148 24464
rect 51188 24424 51189 24464
rect 51147 24415 51189 24424
rect 52107 24464 52149 24473
rect 52107 24424 52108 24464
rect 52148 24424 52149 24464
rect 52107 24415 52149 24424
rect 52587 24464 52629 24473
rect 52587 24424 52588 24464
rect 52628 24424 52629 24464
rect 52587 24415 52629 24424
rect 59107 24464 59165 24465
rect 59107 24424 59116 24464
rect 59156 24424 59165 24464
rect 59107 24423 59165 24424
rect 60843 24464 60885 24473
rect 60843 24424 60844 24464
rect 60884 24424 60885 24464
rect 60843 24415 60885 24424
rect 64779 24464 64821 24473
rect 64779 24424 64780 24464
rect 64820 24424 64821 24464
rect 64779 24415 64821 24424
rect 68523 24464 68565 24473
rect 68523 24424 68524 24464
rect 68564 24424 68565 24464
rect 68523 24415 68565 24424
rect 71211 24464 71253 24473
rect 71211 24424 71212 24464
rect 71252 24424 71253 24464
rect 71211 24415 71253 24424
rect 76099 24464 76157 24465
rect 76099 24424 76108 24464
rect 76148 24424 76157 24464
rect 76099 24423 76157 24424
rect 77163 24464 77205 24473
rect 77163 24424 77164 24464
rect 77204 24424 77205 24464
rect 77163 24415 77205 24424
rect 843 24380 885 24389
rect 843 24340 844 24380
rect 884 24340 885 24380
rect 843 24331 885 24340
rect 32227 24380 32285 24381
rect 32227 24340 32236 24380
rect 32276 24340 32285 24380
rect 32227 24339 32285 24340
rect 39243 24380 39285 24389
rect 39243 24340 39244 24380
rect 39284 24340 39285 24380
rect 39243 24331 39285 24340
rect 40395 24380 40437 24389
rect 40395 24340 40396 24380
rect 40436 24340 40437 24380
rect 40395 24331 40437 24340
rect 44707 24380 44765 24381
rect 44707 24340 44716 24380
rect 44756 24340 44765 24380
rect 44707 24339 44765 24340
rect 50187 24380 50229 24389
rect 50187 24340 50188 24380
rect 50228 24340 50229 24380
rect 50187 24331 50229 24340
rect 50379 24380 50421 24389
rect 50379 24340 50380 24380
rect 50420 24340 50421 24380
rect 50379 24331 50421 24340
rect 576 24212 79584 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 79584 24212
rect 576 24148 79584 24172
rect 2187 24044 2229 24053
rect 2187 24004 2188 24044
rect 2228 24004 2229 24044
rect 2187 23995 2229 24004
rect 35491 24044 35549 24045
rect 35491 24004 35500 24044
rect 35540 24004 35549 24044
rect 35491 24003 35549 24004
rect 35883 24044 35925 24053
rect 35883 24004 35884 24044
rect 35924 24004 35925 24044
rect 35883 23995 35925 24004
rect 43267 24044 43325 24045
rect 43267 24004 43276 24044
rect 43316 24004 43325 24044
rect 43267 24003 43325 24004
rect 44427 24044 44469 24053
rect 44427 24004 44428 24044
rect 44468 24004 44469 24044
rect 44427 23995 44469 24004
rect 55371 24044 55413 24053
rect 55371 24004 55372 24044
rect 55412 24004 55413 24044
rect 55371 23995 55413 24004
rect 28683 23960 28725 23969
rect 28683 23920 28684 23960
rect 28724 23920 28725 23960
rect 28683 23911 28725 23920
rect 32707 23960 32765 23961
rect 32707 23920 32716 23960
rect 32756 23920 32765 23960
rect 32707 23919 32765 23920
rect 37035 23960 37077 23969
rect 37035 23920 37036 23960
rect 37076 23920 37077 23960
rect 37035 23911 37077 23920
rect 45763 23960 45821 23961
rect 45763 23920 45772 23960
rect 45812 23920 45821 23960
rect 45763 23919 45821 23920
rect 46923 23960 46965 23969
rect 46923 23920 46924 23960
rect 46964 23920 46965 23960
rect 46923 23911 46965 23920
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 1795 23876 1853 23877
rect 1795 23836 1804 23876
rect 1844 23836 1853 23876
rect 1795 23835 1853 23836
rect 1987 23876 2045 23877
rect 1987 23836 1996 23876
rect 2036 23836 2045 23876
rect 1987 23835 2045 23836
rect 31459 23876 31517 23877
rect 31459 23836 31468 23876
rect 31508 23836 31517 23876
rect 31459 23835 31517 23836
rect 30699 23792 30741 23801
rect 30699 23752 30700 23792
rect 30740 23752 30741 23792
rect 30699 23743 30741 23752
rect 30891 23792 30933 23801
rect 30891 23752 30892 23792
rect 30932 23752 30933 23792
rect 30891 23743 30933 23752
rect 30979 23792 31037 23793
rect 30979 23752 30988 23792
rect 31028 23752 31037 23792
rect 30979 23751 31037 23752
rect 32035 23792 32093 23793
rect 32035 23752 32044 23792
rect 32084 23752 32093 23792
rect 32035 23751 32093 23752
rect 32331 23792 32373 23801
rect 32331 23752 32332 23792
rect 32372 23752 32373 23792
rect 32331 23743 32373 23752
rect 33475 23792 33533 23793
rect 33475 23752 33484 23792
rect 33524 23752 33533 23792
rect 33475 23751 33533 23752
rect 34339 23792 34397 23793
rect 34339 23752 34348 23792
rect 34388 23752 34397 23792
rect 34339 23751 34397 23752
rect 35883 23792 35925 23801
rect 35883 23752 35884 23792
rect 35924 23752 35925 23792
rect 35883 23743 35925 23752
rect 36075 23792 36117 23801
rect 36075 23752 36076 23792
rect 36116 23752 36117 23792
rect 36075 23743 36117 23752
rect 36163 23792 36221 23793
rect 36163 23752 36172 23792
rect 36212 23752 36221 23792
rect 36163 23751 36221 23752
rect 36355 23792 36413 23793
rect 36355 23752 36364 23792
rect 36404 23752 36413 23792
rect 36355 23751 36413 23752
rect 37315 23792 37373 23793
rect 37315 23752 37324 23792
rect 37364 23752 37373 23792
rect 37315 23751 37373 23752
rect 38859 23792 38901 23801
rect 38859 23752 38860 23792
rect 38900 23752 38901 23792
rect 38859 23743 38901 23752
rect 38955 23792 38997 23801
rect 38955 23752 38956 23792
rect 38996 23752 38997 23792
rect 38955 23743 38997 23752
rect 39051 23792 39093 23801
rect 39051 23752 39052 23792
rect 39092 23752 39093 23792
rect 39051 23743 39093 23752
rect 39339 23792 39381 23801
rect 39339 23752 39340 23792
rect 39380 23752 39381 23792
rect 39339 23743 39381 23752
rect 39531 23792 39573 23801
rect 39531 23752 39532 23792
rect 39572 23752 39573 23792
rect 39531 23743 39573 23752
rect 39619 23792 39677 23793
rect 39619 23752 39628 23792
rect 39668 23752 39677 23792
rect 39619 23751 39677 23752
rect 40483 23792 40541 23793
rect 40483 23752 40492 23792
rect 40532 23752 40541 23792
rect 40483 23751 40541 23752
rect 40683 23792 40725 23801
rect 40683 23752 40684 23792
rect 40724 23752 40725 23792
rect 40683 23743 40725 23752
rect 41251 23792 41309 23793
rect 41251 23752 41260 23792
rect 41300 23752 41309 23792
rect 41251 23751 41309 23752
rect 42115 23792 42173 23793
rect 42115 23752 42124 23792
rect 42164 23752 42173 23792
rect 42115 23751 42173 23752
rect 43947 23792 43989 23801
rect 43947 23752 43948 23792
rect 43988 23752 43989 23792
rect 43947 23743 43989 23752
rect 44043 23792 44085 23801
rect 44043 23752 44044 23792
rect 44084 23752 44085 23792
rect 44043 23743 44085 23752
rect 44139 23792 44181 23801
rect 44139 23752 44140 23792
rect 44180 23752 44181 23792
rect 44139 23743 44181 23752
rect 44235 23792 44277 23801
rect 44235 23752 44236 23792
rect 44276 23752 44277 23792
rect 44235 23743 44277 23752
rect 44427 23792 44469 23801
rect 44427 23752 44428 23792
rect 44468 23752 44469 23792
rect 44427 23743 44469 23752
rect 44619 23792 44661 23801
rect 44619 23752 44620 23792
rect 44660 23752 44661 23792
rect 44619 23743 44661 23752
rect 44707 23792 44765 23793
rect 44707 23752 44716 23792
rect 44756 23752 44765 23792
rect 44707 23751 44765 23752
rect 45091 23792 45149 23793
rect 45091 23752 45100 23792
rect 45140 23752 45149 23792
rect 45091 23751 45149 23752
rect 45387 23792 45429 23801
rect 45387 23752 45388 23792
rect 45428 23752 45429 23792
rect 45387 23743 45429 23752
rect 45483 23792 45525 23801
rect 45483 23752 45484 23792
rect 45524 23752 45525 23792
rect 45483 23743 45525 23752
rect 45963 23792 46005 23801
rect 45963 23752 45964 23792
rect 46004 23752 46005 23792
rect 45963 23743 46005 23752
rect 46059 23792 46101 23801
rect 46059 23752 46060 23792
rect 46100 23752 46101 23792
rect 46059 23743 46101 23752
rect 46147 23792 46205 23793
rect 46147 23752 46156 23792
rect 46196 23752 46205 23792
rect 46147 23751 46205 23752
rect 48355 23792 48413 23793
rect 48355 23752 48364 23792
rect 48404 23752 48413 23792
rect 48355 23751 48413 23752
rect 49219 23792 49277 23793
rect 49219 23752 49228 23792
rect 49268 23752 49277 23792
rect 49219 23751 49277 23752
rect 50571 23792 50613 23801
rect 50571 23752 50572 23792
rect 50612 23752 50613 23792
rect 50571 23743 50613 23752
rect 50763 23792 50805 23801
rect 50763 23752 50764 23792
rect 50804 23752 50805 23792
rect 50763 23743 50805 23752
rect 50851 23792 50909 23793
rect 50851 23752 50860 23792
rect 50900 23752 50909 23792
rect 50851 23751 50909 23752
rect 51051 23792 51093 23801
rect 51051 23752 51052 23792
rect 51092 23752 51093 23792
rect 51051 23743 51093 23752
rect 51243 23792 51285 23801
rect 51243 23752 51244 23792
rect 51284 23752 51285 23792
rect 51243 23743 51285 23752
rect 51331 23792 51389 23793
rect 51331 23752 51340 23792
rect 51380 23752 51389 23792
rect 51331 23751 51389 23752
rect 51723 23792 51765 23801
rect 51723 23752 51724 23792
rect 51764 23752 51765 23792
rect 51723 23743 51765 23752
rect 52099 23792 52157 23793
rect 52099 23752 52108 23792
rect 52148 23752 52157 23792
rect 52099 23751 52157 23752
rect 52963 23792 53021 23793
rect 52963 23752 52972 23792
rect 53012 23752 53021 23792
rect 52963 23751 53021 23752
rect 54787 23792 54845 23793
rect 54787 23752 54796 23792
rect 54836 23752 54845 23792
rect 54787 23751 54845 23752
rect 55075 23792 55133 23793
rect 55075 23752 55084 23792
rect 55124 23752 55133 23792
rect 55075 23751 55133 23752
rect 55371 23792 55413 23801
rect 55371 23752 55372 23792
rect 55412 23752 55413 23792
rect 55371 23743 55413 23752
rect 55563 23792 55605 23801
rect 55563 23752 55564 23792
rect 55604 23752 55605 23792
rect 55563 23743 55605 23752
rect 55651 23792 55709 23793
rect 55651 23752 55660 23792
rect 55700 23752 55709 23792
rect 55651 23751 55709 23752
rect 55843 23792 55901 23793
rect 55843 23752 55852 23792
rect 55892 23752 55901 23792
rect 55843 23751 55901 23752
rect 56131 23792 56189 23793
rect 56131 23752 56140 23792
rect 56180 23752 56189 23792
rect 56131 23751 56189 23752
rect 56419 23792 56477 23793
rect 56419 23752 56428 23792
rect 56468 23752 56477 23792
rect 56419 23751 56477 23752
rect 56803 23792 56861 23793
rect 56803 23752 56812 23792
rect 56852 23752 56861 23792
rect 56803 23751 56861 23752
rect 57283 23792 57341 23793
rect 57283 23752 57292 23792
rect 57332 23752 57341 23792
rect 57283 23751 57341 23752
rect 57667 23792 57725 23793
rect 57667 23752 57676 23792
rect 57716 23752 57725 23792
rect 57667 23751 57725 23752
rect 58051 23792 58109 23793
rect 58051 23752 58060 23792
rect 58100 23752 58109 23792
rect 58051 23751 58109 23752
rect 58435 23792 58493 23793
rect 58435 23752 58444 23792
rect 58484 23752 58493 23792
rect 58435 23751 58493 23752
rect 58915 23792 58973 23793
rect 58915 23752 58924 23792
rect 58964 23752 58973 23792
rect 58915 23751 58973 23752
rect 59299 23792 59357 23793
rect 59299 23752 59308 23792
rect 59348 23752 59357 23792
rect 59299 23751 59357 23752
rect 59683 23792 59741 23793
rect 59683 23752 59692 23792
rect 59732 23752 59741 23792
rect 59683 23751 59741 23752
rect 60067 23792 60125 23793
rect 60067 23752 60076 23792
rect 60116 23752 60125 23792
rect 60067 23751 60125 23752
rect 60451 23792 60509 23793
rect 60451 23752 60460 23792
rect 60500 23752 60509 23792
rect 60451 23751 60509 23752
rect 60835 23792 60893 23793
rect 60835 23752 60844 23792
rect 60884 23752 60893 23792
rect 60835 23751 60893 23752
rect 61315 23792 61373 23793
rect 61315 23752 61324 23792
rect 61364 23752 61373 23792
rect 61315 23751 61373 23752
rect 61699 23792 61757 23793
rect 61699 23752 61708 23792
rect 61748 23752 61757 23792
rect 61699 23751 61757 23752
rect 62083 23792 62141 23793
rect 62083 23752 62092 23792
rect 62132 23752 62141 23792
rect 62083 23751 62141 23752
rect 62467 23792 62525 23793
rect 62467 23752 62476 23792
rect 62516 23752 62525 23792
rect 62467 23751 62525 23752
rect 62851 23792 62909 23793
rect 62851 23752 62860 23792
rect 62900 23752 62909 23792
rect 62851 23751 62909 23752
rect 63235 23792 63293 23793
rect 63235 23752 63244 23792
rect 63284 23752 63293 23792
rect 63235 23751 63293 23752
rect 63715 23792 63773 23793
rect 63715 23752 63724 23792
rect 63764 23752 63773 23792
rect 63715 23751 63773 23752
rect 64099 23792 64157 23793
rect 64099 23752 64108 23792
rect 64148 23752 64157 23792
rect 64099 23751 64157 23752
rect 64483 23792 64541 23793
rect 64483 23752 64492 23792
rect 64532 23752 64541 23792
rect 64483 23751 64541 23752
rect 64867 23792 64925 23793
rect 64867 23752 64876 23792
rect 64916 23752 64925 23792
rect 64867 23751 64925 23752
rect 65251 23792 65309 23793
rect 65251 23752 65260 23792
rect 65300 23752 65309 23792
rect 65251 23751 65309 23752
rect 65731 23792 65789 23793
rect 65731 23752 65740 23792
rect 65780 23752 65789 23792
rect 65731 23751 65789 23752
rect 66115 23792 66173 23793
rect 66115 23752 66124 23792
rect 66164 23752 66173 23792
rect 66115 23751 66173 23752
rect 66499 23792 66557 23793
rect 66499 23752 66508 23792
rect 66548 23752 66557 23792
rect 66499 23751 66557 23752
rect 66883 23792 66941 23793
rect 66883 23752 66892 23792
rect 66932 23752 66941 23792
rect 66883 23751 66941 23752
rect 67267 23792 67325 23793
rect 67267 23752 67276 23792
rect 67316 23752 67325 23792
rect 67267 23751 67325 23752
rect 67747 23792 67805 23793
rect 67747 23752 67756 23792
rect 67796 23752 67805 23792
rect 67747 23751 67805 23752
rect 68131 23792 68189 23793
rect 68131 23752 68140 23792
rect 68180 23752 68189 23792
rect 68131 23751 68189 23752
rect 68515 23792 68573 23793
rect 68515 23752 68524 23792
rect 68564 23752 68573 23792
rect 68515 23751 68573 23752
rect 68899 23792 68957 23793
rect 68899 23752 68908 23792
rect 68948 23752 68957 23792
rect 68899 23751 68957 23752
rect 69283 23792 69341 23793
rect 69283 23752 69292 23792
rect 69332 23752 69341 23792
rect 69283 23751 69341 23752
rect 69763 23792 69821 23793
rect 69763 23752 69772 23792
rect 69812 23752 69821 23792
rect 69763 23751 69821 23752
rect 70147 23792 70205 23793
rect 70147 23752 70156 23792
rect 70196 23752 70205 23792
rect 70147 23751 70205 23752
rect 70531 23792 70589 23793
rect 70531 23752 70540 23792
rect 70580 23752 70589 23792
rect 70531 23751 70589 23752
rect 70915 23792 70973 23793
rect 70915 23752 70924 23792
rect 70964 23752 70973 23792
rect 70915 23751 70973 23752
rect 71299 23792 71357 23793
rect 71299 23752 71308 23792
rect 71348 23752 71357 23792
rect 71299 23751 71357 23752
rect 71683 23792 71741 23793
rect 71683 23752 71692 23792
rect 71732 23752 71741 23792
rect 71683 23751 71741 23752
rect 72067 23792 72125 23793
rect 72067 23752 72076 23792
rect 72116 23752 72125 23792
rect 72067 23751 72125 23752
rect 72451 23792 72509 23793
rect 72451 23752 72460 23792
rect 72500 23752 72509 23792
rect 72451 23751 72509 23752
rect 72835 23792 72893 23793
rect 72835 23752 72844 23792
rect 72884 23752 72893 23792
rect 72835 23751 72893 23752
rect 73315 23792 73373 23793
rect 73315 23752 73324 23792
rect 73364 23752 73373 23792
rect 73315 23751 73373 23752
rect 73699 23792 73757 23793
rect 73699 23752 73708 23792
rect 73748 23752 73757 23792
rect 73699 23751 73757 23752
rect 74083 23792 74141 23793
rect 74083 23752 74092 23792
rect 74132 23752 74141 23792
rect 74083 23751 74141 23752
rect 74467 23792 74525 23793
rect 74467 23752 74476 23792
rect 74516 23752 74525 23792
rect 74467 23751 74525 23752
rect 74851 23792 74909 23793
rect 74851 23752 74860 23792
rect 74900 23752 74909 23792
rect 74851 23751 74909 23752
rect 75235 23792 75293 23793
rect 75235 23752 75244 23792
rect 75284 23752 75293 23792
rect 75235 23751 75293 23752
rect 75619 23792 75677 23793
rect 75619 23752 75628 23792
rect 75668 23752 75677 23792
rect 75619 23751 75677 23752
rect 76099 23792 76157 23793
rect 76099 23752 76108 23792
rect 76148 23752 76157 23792
rect 76099 23751 76157 23752
rect 76963 23792 77021 23793
rect 76963 23752 76972 23792
rect 77012 23752 77021 23792
rect 76963 23751 77021 23752
rect 77251 23792 77309 23793
rect 77251 23752 77260 23792
rect 77300 23752 77309 23792
rect 77251 23751 77309 23752
rect 77443 23792 77501 23793
rect 77443 23752 77452 23792
rect 77492 23752 77501 23792
rect 77443 23751 77501 23752
rect 77731 23792 77789 23793
rect 77731 23752 77740 23792
rect 77780 23752 77789 23792
rect 77731 23751 77789 23752
rect 78115 23792 78173 23793
rect 78115 23752 78124 23792
rect 78164 23752 78173 23792
rect 78115 23751 78173 23752
rect 78499 23792 78557 23793
rect 78499 23752 78508 23792
rect 78548 23752 78557 23792
rect 78499 23751 78557 23752
rect 78787 23792 78845 23793
rect 78787 23752 78796 23792
rect 78836 23752 78845 23792
rect 78787 23751 78845 23752
rect 79075 23792 79133 23793
rect 79075 23752 79084 23792
rect 79124 23752 79133 23792
rect 79075 23751 79133 23752
rect 79363 23792 79421 23793
rect 79363 23752 79372 23792
rect 79412 23752 79421 23792
rect 79363 23751 79421 23752
rect 32427 23708 32469 23717
rect 32427 23668 32428 23708
rect 32468 23668 32469 23708
rect 32427 23659 32469 23668
rect 33099 23708 33141 23717
rect 33099 23668 33100 23708
rect 33140 23668 33141 23708
rect 33099 23659 33141 23668
rect 40587 23708 40629 23717
rect 40587 23668 40588 23708
rect 40628 23668 40629 23708
rect 40587 23659 40629 23668
rect 40875 23708 40917 23717
rect 40875 23668 40876 23708
rect 40916 23668 40917 23708
rect 40875 23659 40917 23668
rect 47979 23708 48021 23717
rect 47979 23668 47980 23708
rect 48020 23668 48021 23708
rect 47979 23659 48021 23668
rect 51147 23708 51189 23717
rect 51147 23668 51148 23708
rect 51188 23668 51189 23708
rect 51147 23659 51189 23668
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 1611 23624 1653 23633
rect 1611 23584 1612 23624
rect 1652 23584 1653 23624
rect 1611 23575 1653 23584
rect 30787 23624 30845 23625
rect 30787 23584 30796 23624
rect 30836 23584 30845 23624
rect 30787 23583 30845 23584
rect 31659 23624 31701 23633
rect 31659 23584 31660 23624
rect 31700 23584 31701 23624
rect 31659 23575 31701 23584
rect 39139 23624 39197 23625
rect 39139 23584 39148 23624
rect 39188 23584 39197 23624
rect 39139 23583 39197 23584
rect 39427 23624 39485 23625
rect 39427 23584 39436 23624
rect 39476 23584 39485 23624
rect 39427 23583 39485 23584
rect 43267 23624 43325 23625
rect 43267 23584 43276 23624
rect 43316 23584 43325 23624
rect 43267 23583 43325 23584
rect 50371 23624 50429 23625
rect 50371 23584 50380 23624
rect 50420 23584 50429 23624
rect 50371 23583 50429 23584
rect 50659 23624 50717 23625
rect 50659 23584 50668 23624
rect 50708 23584 50717 23624
rect 50659 23583 50717 23584
rect 54115 23624 54173 23625
rect 54115 23584 54124 23624
rect 54164 23584 54173 23624
rect 54115 23583 54173 23584
rect 54891 23624 54933 23633
rect 54891 23584 54892 23624
rect 54932 23584 54933 23624
rect 54891 23575 54933 23584
rect 55179 23624 55221 23633
rect 55179 23584 55180 23624
rect 55220 23584 55221 23624
rect 55179 23575 55221 23584
rect 55947 23624 55989 23633
rect 55947 23584 55948 23624
rect 55988 23584 55989 23624
rect 55947 23575 55989 23584
rect 56235 23624 56277 23633
rect 56235 23584 56236 23624
rect 56276 23584 56277 23624
rect 56235 23575 56277 23584
rect 56523 23624 56565 23633
rect 56523 23584 56524 23624
rect 56564 23584 56565 23624
rect 56523 23575 56565 23584
rect 56907 23624 56949 23633
rect 56907 23584 56908 23624
rect 56948 23584 56949 23624
rect 56907 23575 56949 23584
rect 57387 23624 57429 23633
rect 57387 23584 57388 23624
rect 57428 23584 57429 23624
rect 57387 23575 57429 23584
rect 57771 23624 57813 23633
rect 57771 23584 57772 23624
rect 57812 23584 57813 23624
rect 57771 23575 57813 23584
rect 58155 23624 58197 23633
rect 58155 23584 58156 23624
rect 58196 23584 58197 23624
rect 58155 23575 58197 23584
rect 58539 23624 58581 23633
rect 58539 23584 58540 23624
rect 58580 23584 58581 23624
rect 58539 23575 58581 23584
rect 59019 23624 59061 23633
rect 59019 23584 59020 23624
rect 59060 23584 59061 23624
rect 59019 23575 59061 23584
rect 59403 23624 59445 23633
rect 59403 23584 59404 23624
rect 59444 23584 59445 23624
rect 59403 23575 59445 23584
rect 59787 23624 59829 23633
rect 59787 23584 59788 23624
rect 59828 23584 59829 23624
rect 59787 23575 59829 23584
rect 60171 23624 60213 23633
rect 60171 23584 60172 23624
rect 60212 23584 60213 23624
rect 60171 23575 60213 23584
rect 60555 23624 60597 23633
rect 60555 23584 60556 23624
rect 60596 23584 60597 23624
rect 60555 23575 60597 23584
rect 60939 23624 60981 23633
rect 60939 23584 60940 23624
rect 60980 23584 60981 23624
rect 60939 23575 60981 23584
rect 61419 23624 61461 23633
rect 61419 23584 61420 23624
rect 61460 23584 61461 23624
rect 61419 23575 61461 23584
rect 61803 23624 61845 23633
rect 61803 23584 61804 23624
rect 61844 23584 61845 23624
rect 61803 23575 61845 23584
rect 62187 23624 62229 23633
rect 62187 23584 62188 23624
rect 62228 23584 62229 23624
rect 62187 23575 62229 23584
rect 62571 23624 62613 23633
rect 62571 23584 62572 23624
rect 62612 23584 62613 23624
rect 62571 23575 62613 23584
rect 62955 23624 62997 23633
rect 62955 23584 62956 23624
rect 62996 23584 62997 23624
rect 62955 23575 62997 23584
rect 63339 23624 63381 23633
rect 63339 23584 63340 23624
rect 63380 23584 63381 23624
rect 63339 23575 63381 23584
rect 63819 23624 63861 23633
rect 63819 23584 63820 23624
rect 63860 23584 63861 23624
rect 63819 23575 63861 23584
rect 64203 23624 64245 23633
rect 64203 23584 64204 23624
rect 64244 23584 64245 23624
rect 64203 23575 64245 23584
rect 64587 23624 64629 23633
rect 64587 23584 64588 23624
rect 64628 23584 64629 23624
rect 64587 23575 64629 23584
rect 64971 23624 65013 23633
rect 64971 23584 64972 23624
rect 65012 23584 65013 23624
rect 64971 23575 65013 23584
rect 65355 23624 65397 23633
rect 65355 23584 65356 23624
rect 65396 23584 65397 23624
rect 65355 23575 65397 23584
rect 65835 23624 65877 23633
rect 65835 23584 65836 23624
rect 65876 23584 65877 23624
rect 65835 23575 65877 23584
rect 66219 23624 66261 23633
rect 66219 23584 66220 23624
rect 66260 23584 66261 23624
rect 66219 23575 66261 23584
rect 66603 23624 66645 23633
rect 66603 23584 66604 23624
rect 66644 23584 66645 23624
rect 66603 23575 66645 23584
rect 66987 23624 67029 23633
rect 66987 23584 66988 23624
rect 67028 23584 67029 23624
rect 66987 23575 67029 23584
rect 67371 23624 67413 23633
rect 67371 23584 67372 23624
rect 67412 23584 67413 23624
rect 67371 23575 67413 23584
rect 67851 23624 67893 23633
rect 67851 23584 67852 23624
rect 67892 23584 67893 23624
rect 67851 23575 67893 23584
rect 68235 23624 68277 23633
rect 68235 23584 68236 23624
rect 68276 23584 68277 23624
rect 68235 23575 68277 23584
rect 68619 23624 68661 23633
rect 68619 23584 68620 23624
rect 68660 23584 68661 23624
rect 68619 23575 68661 23584
rect 69003 23624 69045 23633
rect 69003 23584 69004 23624
rect 69044 23584 69045 23624
rect 69003 23575 69045 23584
rect 69387 23624 69429 23633
rect 69387 23584 69388 23624
rect 69428 23584 69429 23624
rect 69387 23575 69429 23584
rect 69867 23624 69909 23633
rect 69867 23584 69868 23624
rect 69908 23584 69909 23624
rect 69867 23575 69909 23584
rect 70251 23624 70293 23633
rect 70251 23584 70252 23624
rect 70292 23584 70293 23624
rect 70251 23575 70293 23584
rect 70635 23624 70677 23633
rect 70635 23584 70636 23624
rect 70676 23584 70677 23624
rect 70635 23575 70677 23584
rect 71019 23624 71061 23633
rect 71019 23584 71020 23624
rect 71060 23584 71061 23624
rect 71019 23575 71061 23584
rect 71403 23624 71445 23633
rect 71403 23584 71404 23624
rect 71444 23584 71445 23624
rect 71403 23575 71445 23584
rect 71787 23624 71829 23633
rect 71787 23584 71788 23624
rect 71828 23584 71829 23624
rect 71787 23575 71829 23584
rect 72171 23624 72213 23633
rect 72171 23584 72172 23624
rect 72212 23584 72213 23624
rect 72171 23575 72213 23584
rect 72555 23624 72597 23633
rect 72555 23584 72556 23624
rect 72596 23584 72597 23624
rect 72555 23575 72597 23584
rect 72939 23624 72981 23633
rect 72939 23584 72940 23624
rect 72980 23584 72981 23624
rect 72939 23575 72981 23584
rect 73419 23624 73461 23633
rect 73419 23584 73420 23624
rect 73460 23584 73461 23624
rect 73419 23575 73461 23584
rect 73803 23624 73845 23633
rect 73803 23584 73804 23624
rect 73844 23584 73845 23624
rect 73803 23575 73845 23584
rect 74187 23624 74229 23633
rect 74187 23584 74188 23624
rect 74228 23584 74229 23624
rect 74187 23575 74229 23584
rect 74571 23624 74613 23633
rect 74571 23584 74572 23624
rect 74612 23584 74613 23624
rect 74571 23575 74613 23584
rect 74955 23624 74997 23633
rect 74955 23584 74956 23624
rect 74996 23584 74997 23624
rect 74955 23575 74997 23584
rect 75339 23624 75381 23633
rect 75339 23584 75340 23624
rect 75380 23584 75381 23624
rect 75339 23575 75381 23584
rect 75723 23624 75765 23633
rect 75723 23584 75724 23624
rect 75764 23584 75765 23624
rect 75723 23575 75765 23584
rect 76203 23624 76245 23633
rect 76203 23584 76204 23624
rect 76244 23584 76245 23624
rect 76203 23575 76245 23584
rect 76875 23624 76917 23633
rect 76875 23584 76876 23624
rect 76916 23584 76917 23624
rect 76875 23575 76917 23584
rect 77163 23624 77205 23633
rect 77163 23584 77164 23624
rect 77204 23584 77205 23624
rect 77163 23575 77205 23584
rect 77547 23624 77589 23633
rect 77547 23584 77548 23624
rect 77588 23584 77589 23624
rect 77547 23575 77589 23584
rect 77835 23624 77877 23633
rect 77835 23584 77836 23624
rect 77876 23584 77877 23624
rect 77835 23575 77877 23584
rect 78219 23624 78261 23633
rect 78219 23584 78220 23624
rect 78260 23584 78261 23624
rect 78219 23575 78261 23584
rect 78603 23624 78645 23633
rect 78603 23584 78604 23624
rect 78644 23584 78645 23624
rect 78603 23575 78645 23584
rect 78891 23624 78933 23633
rect 78891 23584 78892 23624
rect 78932 23584 78933 23624
rect 78891 23575 78933 23584
rect 79179 23624 79221 23633
rect 79179 23584 79180 23624
rect 79220 23584 79221 23624
rect 79179 23575 79221 23584
rect 79467 23624 79509 23633
rect 79467 23584 79468 23624
rect 79508 23584 79509 23624
rect 79467 23575 79509 23584
rect 576 23456 79584 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 79584 23456
rect 576 23392 79584 23416
rect 41067 23330 41109 23339
rect 41067 23290 41068 23330
rect 41108 23290 41109 23330
rect 31267 23288 31325 23289
rect 31267 23248 31276 23288
rect 31316 23248 31325 23288
rect 31267 23247 31325 23248
rect 32803 23288 32861 23289
rect 32803 23248 32812 23288
rect 32852 23248 32861 23288
rect 32803 23247 32861 23248
rect 35683 23288 35741 23289
rect 35683 23248 35692 23288
rect 35732 23248 35741 23288
rect 35683 23247 35741 23248
rect 37891 23288 37949 23289
rect 37891 23248 37900 23288
rect 37940 23248 37949 23288
rect 37891 23247 37949 23248
rect 40867 23288 40925 23289
rect 40867 23248 40876 23288
rect 40916 23248 40925 23288
rect 41067 23281 41109 23290
rect 44707 23288 44765 23289
rect 40867 23247 40925 23248
rect 44707 23248 44716 23288
rect 44756 23248 44765 23288
rect 44707 23247 44765 23248
rect 48835 23288 48893 23289
rect 48835 23248 48844 23288
rect 48884 23248 48893 23288
rect 48835 23247 48893 23248
rect 49515 23288 49557 23297
rect 49515 23248 49516 23288
rect 49556 23248 49557 23288
rect 49515 23239 49557 23248
rect 49987 23288 50045 23289
rect 49987 23248 49996 23288
rect 50036 23248 50045 23288
rect 49987 23247 50045 23248
rect 28203 23204 28245 23213
rect 28203 23164 28204 23204
rect 28244 23164 28245 23204
rect 28203 23155 28245 23164
rect 32427 23204 32469 23213
rect 32427 23164 32428 23204
rect 32468 23164 32469 23204
rect 32427 23155 32469 23164
rect 36651 23204 36693 23213
rect 36651 23164 36652 23204
rect 36692 23164 36693 23204
rect 36651 23155 36693 23164
rect 37227 23204 37269 23213
rect 37227 23164 37228 23204
rect 37268 23164 37269 23204
rect 37227 23155 37269 23164
rect 41355 23204 41397 23213
rect 41355 23164 41356 23204
rect 41396 23164 41397 23204
rect 41355 23155 41397 23164
rect 50667 23204 50709 23213
rect 50667 23164 50668 23204
rect 50708 23164 50709 23204
rect 50667 23155 50709 23164
rect 51243 23204 51285 23213
rect 51243 23164 51244 23204
rect 51284 23164 51285 23204
rect 51243 23155 51285 23164
rect 51627 23204 51669 23213
rect 51627 23164 51628 23204
rect 51668 23164 51669 23204
rect 51627 23155 51669 23164
rect 51523 23141 51581 23142
rect 1515 23120 1557 23129
rect 1515 23080 1516 23120
rect 1556 23080 1557 23120
rect 1515 23071 1557 23080
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 1941 23120
rect 1899 23071 1941 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 28579 23120 28637 23121
rect 28579 23080 28588 23120
rect 28628 23080 28637 23120
rect 28579 23079 28637 23080
rect 29443 23120 29501 23121
rect 29443 23080 29452 23120
rect 29492 23080 29501 23120
rect 29443 23079 29501 23080
rect 31179 23120 31221 23129
rect 31179 23080 31180 23120
rect 31220 23080 31221 23120
rect 31179 23071 31221 23080
rect 31371 23120 31413 23129
rect 31371 23080 31372 23120
rect 31412 23080 31413 23120
rect 31371 23071 31413 23080
rect 31459 23120 31517 23121
rect 31459 23080 31468 23120
rect 31508 23080 31517 23120
rect 31459 23079 31517 23080
rect 32323 23120 32381 23121
rect 32323 23080 32332 23120
rect 32372 23080 32381 23120
rect 32323 23079 32381 23080
rect 32523 23120 32565 23129
rect 32523 23080 32524 23120
rect 32564 23080 32565 23120
rect 32523 23071 32565 23080
rect 32715 23120 32757 23129
rect 32715 23080 32716 23120
rect 32756 23080 32757 23120
rect 32715 23071 32757 23080
rect 32907 23120 32949 23129
rect 32907 23080 32908 23120
rect 32948 23080 32949 23120
rect 32907 23071 32949 23080
rect 32995 23120 33053 23121
rect 32995 23080 33004 23120
rect 33044 23080 33053 23120
rect 32995 23079 33053 23080
rect 33187 23120 33245 23121
rect 33187 23080 33196 23120
rect 33236 23080 33245 23120
rect 33187 23079 33245 23080
rect 33291 23120 33333 23129
rect 33291 23080 33292 23120
rect 33332 23080 33333 23120
rect 33291 23071 33333 23080
rect 33387 23120 33429 23129
rect 33387 23080 33388 23120
rect 33428 23080 33429 23120
rect 33387 23071 33429 23080
rect 35787 23120 35829 23129
rect 35787 23080 35788 23120
rect 35828 23080 35829 23120
rect 35787 23071 35829 23080
rect 35883 23120 35925 23129
rect 35883 23080 35884 23120
rect 35924 23080 35925 23120
rect 35883 23071 35925 23080
rect 35979 23120 36021 23129
rect 35979 23080 35980 23120
rect 36020 23080 36021 23120
rect 35979 23071 36021 23080
rect 36259 23120 36317 23121
rect 36259 23080 36268 23120
rect 36308 23080 36317 23120
rect 36259 23079 36317 23080
rect 36555 23120 36597 23129
rect 36555 23080 36556 23120
rect 36596 23080 36597 23120
rect 36555 23071 36597 23080
rect 37131 23120 37173 23129
rect 37131 23080 37132 23120
rect 37172 23080 37173 23120
rect 37131 23071 37173 23080
rect 37315 23120 37373 23121
rect 37315 23080 37324 23120
rect 37364 23080 37373 23120
rect 37315 23079 37373 23080
rect 37803 23120 37845 23129
rect 37803 23080 37804 23120
rect 37844 23080 37845 23120
rect 37803 23071 37845 23080
rect 37995 23120 38037 23129
rect 37995 23080 37996 23120
rect 38036 23080 38037 23120
rect 37995 23071 38037 23080
rect 38083 23120 38141 23121
rect 38083 23080 38092 23120
rect 38132 23080 38141 23120
rect 38083 23079 38141 23080
rect 38475 23120 38517 23129
rect 38475 23080 38476 23120
rect 38516 23080 38517 23120
rect 38475 23071 38517 23080
rect 38851 23120 38909 23121
rect 38851 23080 38860 23120
rect 38900 23080 38909 23120
rect 38851 23079 38909 23080
rect 39715 23120 39773 23121
rect 39715 23080 39724 23120
rect 39764 23080 39773 23120
rect 39715 23079 39773 23080
rect 41451 23120 41493 23129
rect 41451 23080 41452 23120
rect 41492 23080 41493 23120
rect 41451 23071 41493 23080
rect 41731 23120 41789 23121
rect 41731 23080 41740 23120
rect 41780 23080 41789 23120
rect 41731 23079 41789 23080
rect 44619 23120 44661 23129
rect 44619 23080 44620 23120
rect 44660 23080 44661 23120
rect 44619 23071 44661 23080
rect 44811 23120 44853 23129
rect 44811 23080 44812 23120
rect 44852 23080 44853 23120
rect 44811 23071 44853 23080
rect 44899 23120 44957 23121
rect 44899 23080 44908 23120
rect 44948 23080 44957 23120
rect 44899 23079 44957 23080
rect 45483 23120 45525 23129
rect 45483 23080 45484 23120
rect 45524 23080 45525 23120
rect 45483 23071 45525 23080
rect 45579 23120 45621 23129
rect 45579 23080 45580 23120
rect 45620 23080 45621 23120
rect 45579 23071 45621 23080
rect 45667 23120 45725 23121
rect 45667 23080 45676 23120
rect 45716 23080 45725 23120
rect 45667 23079 45725 23080
rect 45859 23120 45917 23121
rect 45859 23080 45868 23120
rect 45908 23080 45917 23120
rect 45859 23079 45917 23080
rect 45963 23120 46005 23129
rect 45963 23080 45964 23120
rect 46004 23080 46005 23120
rect 46443 23120 46485 23129
rect 45963 23071 46005 23080
rect 46155 23109 46197 23118
rect 46155 23069 46156 23109
rect 46196 23069 46197 23109
rect 46443 23080 46444 23120
rect 46484 23080 46485 23120
rect 46443 23071 46485 23080
rect 46819 23120 46877 23121
rect 46819 23080 46828 23120
rect 46868 23080 46877 23120
rect 46819 23079 46877 23080
rect 47683 23120 47741 23121
rect 47683 23080 47692 23120
rect 47732 23080 47741 23120
rect 47683 23079 47741 23080
rect 49707 23120 49749 23129
rect 49707 23080 49708 23120
rect 49748 23080 49749 23120
rect 49707 23071 49749 23080
rect 49803 23120 49845 23129
rect 49803 23080 49804 23120
rect 49844 23080 49845 23120
rect 49803 23071 49845 23080
rect 49899 23120 49941 23129
rect 49899 23080 49900 23120
rect 49940 23080 49941 23120
rect 49899 23071 49941 23080
rect 50275 23120 50333 23121
rect 50275 23080 50284 23120
rect 50324 23080 50333 23120
rect 50275 23079 50333 23080
rect 50571 23120 50613 23129
rect 50571 23080 50572 23120
rect 50612 23080 50613 23120
rect 50571 23071 50613 23080
rect 51147 23120 51189 23129
rect 51147 23080 51148 23120
rect 51188 23080 51189 23120
rect 51147 23071 51189 23080
rect 51331 23120 51389 23121
rect 51331 23080 51340 23120
rect 51380 23080 51389 23120
rect 51523 23101 51532 23141
rect 51572 23101 51581 23141
rect 51523 23100 51581 23101
rect 51723 23120 51765 23129
rect 51331 23079 51389 23080
rect 51723 23080 51724 23120
rect 51764 23080 51765 23120
rect 51723 23071 51765 23080
rect 52579 23120 52637 23121
rect 52579 23080 52588 23120
rect 52628 23080 52637 23120
rect 52579 23079 52637 23080
rect 52683 23120 52725 23129
rect 52683 23080 52684 23120
rect 52724 23080 52725 23120
rect 52683 23071 52725 23080
rect 46155 23060 46197 23069
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 42403 23036 42461 23037
rect 42403 22996 42412 23036
rect 42452 22996 42461 23036
rect 42403 22995 42461 22996
rect 49315 23036 49373 23037
rect 49315 22996 49324 23036
rect 49364 22996 49373 23036
rect 49315 22995 49373 22996
rect 1515 22952 1557 22961
rect 1515 22912 1516 22952
rect 1556 22912 1557 22952
rect 1515 22903 1557 22912
rect 33579 22952 33621 22961
rect 33579 22912 33580 22952
rect 33620 22912 33621 22952
rect 33579 22903 33621 22912
rect 35499 22952 35541 22961
rect 35499 22912 35500 22952
rect 35540 22912 35541 22952
rect 35499 22903 35541 22912
rect 36931 22952 36989 22953
rect 36931 22912 36940 22952
rect 36980 22912 36989 22952
rect 36931 22911 36989 22912
rect 42027 22952 42069 22961
rect 42027 22912 42028 22952
rect 42068 22912 42069 22952
rect 42027 22903 42069 22912
rect 42795 22952 42837 22961
rect 42795 22912 42796 22952
rect 42836 22912 42837 22952
rect 42795 22903 42837 22912
rect 50947 22952 51005 22953
rect 50947 22912 50956 22952
rect 50996 22912 51005 22952
rect 50947 22911 51005 22912
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 1707 22868 1749 22877
rect 1707 22828 1708 22868
rect 1748 22828 1749 22868
rect 1707 22819 1749 22828
rect 1899 22868 1941 22877
rect 1899 22828 1900 22868
rect 1940 22828 1941 22868
rect 1899 22819 1941 22828
rect 30595 22868 30653 22869
rect 30595 22828 30604 22868
rect 30644 22828 30653 22868
rect 30595 22827 30653 22828
rect 42603 22868 42645 22877
rect 42603 22828 42604 22868
rect 42644 22828 42645 22868
rect 42603 22819 42645 22828
rect 46155 22868 46197 22877
rect 46155 22828 46156 22868
rect 46196 22828 46197 22868
rect 46155 22819 46197 22828
rect 49515 22868 49557 22877
rect 49515 22828 49516 22868
rect 49556 22828 49557 22868
rect 49515 22819 49557 22828
rect 576 22700 52800 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 52800 22700
rect 576 22636 52800 22660
rect 34915 22532 34973 22533
rect 34915 22492 34924 22532
rect 34964 22492 34973 22532
rect 34915 22491 34973 22492
rect 39051 22532 39093 22541
rect 39051 22492 39052 22532
rect 39092 22492 39093 22532
rect 39051 22483 39093 22492
rect 43459 22532 43517 22533
rect 43459 22492 43468 22532
rect 43508 22492 43517 22532
rect 43459 22491 43517 22492
rect 51243 22532 51285 22541
rect 51243 22492 51244 22532
rect 51284 22492 51285 22532
rect 51243 22483 51285 22492
rect 52011 22532 52053 22541
rect 52011 22492 52012 22532
rect 52052 22492 52053 22532
rect 52011 22483 52053 22492
rect 52395 22532 52437 22541
rect 52395 22492 52396 22532
rect 52436 22492 52437 22532
rect 52395 22483 52437 22492
rect 52683 22532 52725 22541
rect 52683 22492 52684 22532
rect 52724 22492 52725 22532
rect 52683 22483 52725 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 31555 22448 31613 22449
rect 31555 22408 31564 22448
rect 31604 22408 31613 22448
rect 31555 22407 31613 22408
rect 35595 22448 35637 22457
rect 35595 22408 35596 22448
rect 35636 22408 35637 22448
rect 35595 22399 35637 22408
rect 38179 22448 38237 22449
rect 38179 22408 38188 22448
rect 38228 22408 38237 22448
rect 38179 22407 38237 22408
rect 38859 22448 38901 22457
rect 38859 22408 38860 22448
rect 38900 22408 38901 22448
rect 38859 22399 38901 22408
rect 40395 22448 40437 22457
rect 40395 22408 40396 22448
rect 40436 22408 40437 22448
rect 40395 22399 40437 22408
rect 46443 22448 46485 22457
rect 46443 22408 46444 22448
rect 46484 22408 46485 22448
rect 46443 22399 46485 22408
rect 48171 22448 48213 22457
rect 48171 22408 48172 22448
rect 48212 22408 48213 22448
rect 48171 22399 48213 22408
rect 3235 22364 3293 22365
rect 3235 22324 3244 22364
rect 3284 22324 3293 22364
rect 3235 22323 3293 22324
rect 28003 22364 28061 22365
rect 28003 22324 28012 22364
rect 28052 22324 28061 22364
rect 28003 22323 28061 22324
rect 40195 22364 40253 22365
rect 40195 22324 40204 22364
rect 40244 22324 40253 22364
rect 40195 22323 40253 22324
rect 49027 22364 49085 22365
rect 49027 22324 49036 22364
rect 49076 22324 49085 22364
rect 49027 22323 49085 22324
rect 30315 22280 30357 22289
rect 30315 22240 30316 22280
rect 30356 22240 30357 22280
rect 30315 22231 30357 22240
rect 30411 22280 30453 22289
rect 30411 22240 30412 22280
rect 30452 22240 30453 22280
rect 30411 22231 30453 22240
rect 30507 22280 30549 22289
rect 30507 22240 30508 22280
rect 30548 22240 30549 22280
rect 30507 22231 30549 22240
rect 30603 22280 30645 22289
rect 30603 22240 30604 22280
rect 30644 22240 30645 22280
rect 30603 22231 30645 22240
rect 30883 22280 30941 22281
rect 30883 22240 30892 22280
rect 30932 22240 30941 22280
rect 30883 22239 30941 22240
rect 31179 22280 31221 22289
rect 31179 22240 31180 22280
rect 31220 22240 31221 22280
rect 31179 22231 31221 22240
rect 31275 22280 31317 22289
rect 31275 22240 31276 22280
rect 31316 22240 31317 22280
rect 31275 22231 31317 22240
rect 31851 22280 31893 22289
rect 31851 22240 31852 22280
rect 31892 22240 31893 22280
rect 31851 22231 31893 22240
rect 32043 22280 32085 22289
rect 32043 22240 32044 22280
rect 32084 22240 32085 22280
rect 32043 22231 32085 22240
rect 32131 22280 32189 22281
rect 32131 22240 32140 22280
rect 32180 22240 32189 22280
rect 32131 22239 32189 22240
rect 32899 22280 32957 22281
rect 32899 22240 32908 22280
rect 32948 22240 32957 22280
rect 32899 22239 32957 22240
rect 33763 22280 33821 22281
rect 33763 22240 33772 22280
rect 33812 22240 33821 22280
rect 33763 22239 33821 22240
rect 36163 22280 36221 22281
rect 36163 22240 36172 22280
rect 36212 22240 36221 22280
rect 36163 22239 36221 22240
rect 37027 22280 37085 22281
rect 37027 22240 37036 22280
rect 37076 22240 37085 22280
rect 37027 22239 37085 22240
rect 39051 22280 39093 22289
rect 39051 22240 39052 22280
rect 39092 22240 39093 22280
rect 39051 22231 39093 22240
rect 39243 22280 39285 22289
rect 39243 22240 39244 22280
rect 39284 22240 39285 22280
rect 39243 22231 39285 22240
rect 39331 22280 39389 22281
rect 39331 22240 39340 22280
rect 39380 22240 39389 22280
rect 39331 22239 39389 22240
rect 40587 22280 40629 22289
rect 40587 22240 40588 22280
rect 40628 22240 40629 22280
rect 40587 22231 40629 22240
rect 40779 22280 40821 22289
rect 40779 22240 40780 22280
rect 40820 22240 40821 22280
rect 40779 22231 40821 22240
rect 40867 22280 40925 22281
rect 40867 22240 40876 22280
rect 40916 22240 40925 22280
rect 40867 22239 40925 22240
rect 41443 22280 41501 22281
rect 41443 22240 41452 22280
rect 41492 22240 41501 22280
rect 41443 22239 41501 22240
rect 42307 22280 42365 22281
rect 42307 22240 42316 22280
rect 42356 22240 42365 22280
rect 42307 22239 42365 22240
rect 45099 22280 45141 22289
rect 45099 22240 45100 22280
rect 45140 22240 45141 22280
rect 45099 22231 45141 22240
rect 45291 22280 45333 22289
rect 45291 22240 45292 22280
rect 45332 22240 45333 22280
rect 45291 22231 45333 22240
rect 45379 22280 45437 22281
rect 45379 22240 45388 22280
rect 45428 22240 45437 22280
rect 45379 22239 45437 22240
rect 45579 22280 45621 22289
rect 45579 22240 45580 22280
rect 45620 22240 45621 22280
rect 45579 22231 45621 22240
rect 45763 22280 45821 22281
rect 45763 22240 45772 22280
rect 45812 22240 45821 22280
rect 45763 22239 45821 22240
rect 48555 22280 48597 22289
rect 48555 22240 48556 22280
rect 48596 22240 48597 22280
rect 48555 22231 48597 22240
rect 48651 22280 48693 22289
rect 48651 22240 48652 22280
rect 48692 22240 48693 22280
rect 48651 22231 48693 22240
rect 48747 22280 48789 22289
rect 48747 22240 48748 22280
rect 48788 22240 48789 22280
rect 48747 22231 48789 22240
rect 49419 22280 49461 22289
rect 49419 22240 49420 22280
rect 49460 22240 49461 22280
rect 49419 22231 49461 22240
rect 49611 22280 49653 22289
rect 49611 22240 49612 22280
rect 49652 22240 49653 22280
rect 49611 22231 49653 22240
rect 49699 22280 49757 22281
rect 49699 22240 49708 22280
rect 49748 22240 49757 22280
rect 49699 22239 49757 22240
rect 50179 22280 50237 22281
rect 50179 22240 50188 22280
rect 50228 22240 50237 22280
rect 50179 22239 50237 22240
rect 50379 22280 50421 22289
rect 50379 22240 50380 22280
rect 50420 22240 50421 22280
rect 50379 22231 50421 22240
rect 51435 22280 51477 22289
rect 51435 22240 51436 22280
rect 51476 22240 51477 22280
rect 51435 22231 51477 22240
rect 52099 22280 52157 22281
rect 52099 22240 52108 22280
rect 52148 22240 52157 22280
rect 52099 22239 52157 22240
rect 52291 22280 52349 22281
rect 52291 22240 52300 22280
rect 52340 22240 52349 22280
rect 52291 22239 52349 22240
rect 52579 22280 52637 22281
rect 52579 22240 52588 22280
rect 52628 22240 52637 22280
rect 52579 22239 52637 22240
rect 32523 22196 32565 22205
rect 32523 22156 32524 22196
rect 32564 22156 32565 22196
rect 32523 22147 32565 22156
rect 35787 22196 35829 22205
rect 35787 22156 35788 22196
rect 35828 22156 35829 22196
rect 35787 22147 35829 22156
rect 41067 22196 41109 22205
rect 41067 22156 41068 22196
rect 41108 22156 41109 22196
rect 41067 22147 41109 22156
rect 45675 22196 45717 22205
rect 45675 22156 45676 22196
rect 45716 22156 45717 22196
rect 45675 22147 45717 22156
rect 50283 22196 50325 22205
rect 50283 22156 50284 22196
rect 50324 22156 50325 22196
rect 50283 22147 50325 22156
rect 3435 22112 3477 22121
rect 3435 22072 3436 22112
rect 3476 22072 3477 22112
rect 3435 22063 3477 22072
rect 28203 22112 28245 22121
rect 28203 22072 28204 22112
rect 28244 22072 28245 22112
rect 28203 22063 28245 22072
rect 31939 22112 31997 22113
rect 31939 22072 31948 22112
rect 31988 22072 31997 22112
rect 31939 22071 31997 22072
rect 34915 22112 34973 22113
rect 34915 22072 34924 22112
rect 34964 22072 34973 22112
rect 34915 22071 34973 22072
rect 40675 22112 40733 22113
rect 40675 22072 40684 22112
rect 40724 22072 40733 22112
rect 40675 22071 40733 22072
rect 45187 22112 45245 22113
rect 45187 22072 45196 22112
rect 45236 22072 45245 22112
rect 45187 22071 45245 22072
rect 48835 22112 48893 22113
rect 48835 22072 48844 22112
rect 48884 22072 48893 22112
rect 48835 22071 48893 22072
rect 49227 22112 49269 22121
rect 49227 22072 49228 22112
rect 49268 22072 49269 22112
rect 49227 22063 49269 22072
rect 49507 22112 49565 22113
rect 49507 22072 49516 22112
rect 49556 22072 49565 22112
rect 49507 22071 49565 22072
rect 576 21944 52800 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 52800 21944
rect 576 21880 52800 21904
rect 3235 21776 3293 21777
rect 3235 21736 3244 21776
rect 3284 21736 3293 21776
rect 3235 21735 3293 21736
rect 29443 21776 29501 21777
rect 29443 21736 29452 21776
rect 29492 21736 29501 21776
rect 29443 21735 29501 21736
rect 36259 21776 36317 21777
rect 36259 21736 36268 21776
rect 36308 21736 36317 21776
rect 36259 21735 36317 21736
rect 44707 21776 44765 21777
rect 44707 21736 44716 21776
rect 44756 21736 44765 21776
rect 44707 21735 44765 21736
rect 31563 21692 31605 21701
rect 31563 21652 31564 21692
rect 31604 21652 31605 21692
rect 31563 21643 31605 21652
rect 32139 21692 32181 21701
rect 32139 21652 32140 21692
rect 32180 21652 32181 21692
rect 32139 21643 32181 21652
rect 41163 21692 41205 21701
rect 41163 21652 41164 21692
rect 41204 21652 41205 21692
rect 41163 21643 41205 21652
rect 42315 21692 42357 21701
rect 42315 21652 42316 21692
rect 42356 21652 42357 21692
rect 42315 21643 42357 21652
rect 51051 21692 51093 21701
rect 51051 21652 51052 21692
rect 51092 21652 51093 21692
rect 51051 21643 51093 21652
rect 3043 21608 3101 21609
rect 3043 21568 3052 21608
rect 3092 21568 3101 21608
rect 3043 21567 3101 21568
rect 3147 21608 3189 21617
rect 3147 21568 3148 21608
rect 3188 21568 3189 21608
rect 3147 21559 3189 21568
rect 3339 21608 3381 21617
rect 3339 21568 3340 21608
rect 3380 21568 3381 21608
rect 3339 21559 3381 21568
rect 27819 21608 27861 21617
rect 27819 21568 27820 21608
rect 27860 21568 27861 21608
rect 27819 21559 27861 21568
rect 27915 21608 27957 21617
rect 27915 21568 27916 21608
rect 27956 21568 27957 21608
rect 27915 21559 27957 21568
rect 28011 21608 28053 21617
rect 28011 21568 28012 21608
rect 28052 21568 28053 21608
rect 28011 21559 28053 21568
rect 28107 21608 28149 21617
rect 28107 21568 28108 21608
rect 28148 21568 28149 21608
rect 28107 21559 28149 21568
rect 28299 21608 28341 21617
rect 28299 21568 28300 21608
rect 28340 21568 28341 21608
rect 28299 21559 28341 21568
rect 28491 21608 28533 21617
rect 28491 21568 28492 21608
rect 28532 21568 28533 21608
rect 28491 21559 28533 21568
rect 28579 21608 28637 21609
rect 28579 21568 28588 21608
rect 28628 21568 28637 21608
rect 28579 21567 28637 21568
rect 28875 21608 28917 21617
rect 28875 21568 28876 21608
rect 28916 21568 28917 21608
rect 28875 21559 28917 21568
rect 29059 21608 29117 21609
rect 29059 21568 29068 21608
rect 29108 21568 29117 21608
rect 29059 21567 29117 21568
rect 29355 21608 29397 21617
rect 29355 21568 29356 21608
rect 29396 21568 29397 21608
rect 29355 21559 29397 21568
rect 29547 21608 29589 21617
rect 29547 21568 29548 21608
rect 29588 21568 29589 21608
rect 29547 21559 29589 21568
rect 29635 21608 29693 21609
rect 29635 21568 29644 21608
rect 29684 21568 29693 21608
rect 29635 21567 29693 21568
rect 31459 21608 31517 21609
rect 31459 21568 31468 21608
rect 31508 21568 31517 21608
rect 31459 21567 31517 21568
rect 31659 21608 31701 21617
rect 31659 21568 31660 21608
rect 31700 21568 31701 21608
rect 31659 21559 31701 21568
rect 32043 21608 32085 21617
rect 32043 21568 32044 21608
rect 32084 21568 32085 21608
rect 32043 21559 32085 21568
rect 32227 21608 32285 21609
rect 32227 21568 32236 21608
rect 32276 21568 32285 21608
rect 32227 21567 32285 21568
rect 36171 21608 36213 21617
rect 36171 21568 36172 21608
rect 36212 21568 36213 21608
rect 36171 21559 36213 21568
rect 36363 21608 36405 21617
rect 36363 21568 36364 21608
rect 36404 21568 36405 21608
rect 36363 21559 36405 21568
rect 36451 21608 36509 21609
rect 36451 21568 36460 21608
rect 36500 21568 36509 21608
rect 36451 21567 36509 21568
rect 36643 21608 36701 21609
rect 36643 21568 36652 21608
rect 36692 21568 36701 21608
rect 36643 21567 36701 21568
rect 36843 21608 36885 21617
rect 36843 21568 36844 21608
rect 36884 21568 36885 21608
rect 36843 21559 36885 21568
rect 39051 21608 39093 21617
rect 39051 21568 39052 21608
rect 39092 21568 39093 21608
rect 39051 21559 39093 21568
rect 39147 21608 39189 21617
rect 39147 21568 39148 21608
rect 39188 21568 39189 21608
rect 39147 21559 39189 21568
rect 39243 21608 39285 21617
rect 39243 21568 39244 21608
rect 39284 21568 39285 21608
rect 39243 21559 39285 21568
rect 39339 21608 39381 21617
rect 39339 21568 39340 21608
rect 39380 21568 39381 21608
rect 39339 21559 39381 21568
rect 41059 21608 41117 21609
rect 41059 21568 41068 21608
rect 41108 21568 41117 21608
rect 41059 21567 41117 21568
rect 41259 21608 41301 21617
rect 41259 21568 41260 21608
rect 41300 21568 41301 21608
rect 41259 21559 41301 21568
rect 42691 21608 42749 21609
rect 42691 21568 42700 21608
rect 42740 21568 42749 21608
rect 42691 21567 42749 21568
rect 43555 21608 43613 21609
rect 43555 21568 43564 21608
rect 43604 21568 43613 21608
rect 43555 21567 43613 21568
rect 44995 21608 45053 21609
rect 44995 21568 45004 21608
rect 45044 21568 45053 21608
rect 44995 21567 45053 21568
rect 45291 21608 45333 21617
rect 45291 21568 45292 21608
rect 45332 21568 45333 21608
rect 45291 21559 45333 21568
rect 45387 21608 45429 21617
rect 45387 21568 45388 21608
rect 45428 21568 45429 21608
rect 45387 21559 45429 21568
rect 45963 21608 46005 21617
rect 45963 21568 45964 21608
rect 46004 21568 46005 21608
rect 45963 21559 46005 21568
rect 46339 21608 46397 21609
rect 46339 21568 46348 21608
rect 46388 21568 46397 21608
rect 46339 21567 46397 21568
rect 47203 21608 47261 21609
rect 47203 21568 47212 21608
rect 47252 21568 47261 21608
rect 47203 21567 47261 21568
rect 48843 21608 48885 21617
rect 48843 21568 48844 21608
rect 48884 21568 48885 21608
rect 48843 21559 48885 21568
rect 49035 21608 49077 21617
rect 49035 21568 49036 21608
rect 49076 21568 49077 21608
rect 49035 21559 49077 21568
rect 49123 21608 49181 21609
rect 49123 21568 49132 21608
rect 49172 21568 49181 21608
rect 49123 21567 49181 21568
rect 49507 21608 49565 21609
rect 49507 21568 49516 21608
rect 49556 21568 49565 21608
rect 49507 21567 49565 21568
rect 49611 21608 49653 21617
rect 49611 21568 49612 21608
rect 49652 21568 49653 21608
rect 49611 21559 49653 21568
rect 49707 21608 49749 21617
rect 49707 21568 49708 21608
rect 49748 21568 49749 21608
rect 49707 21559 49749 21568
rect 50187 21608 50229 21617
rect 50187 21568 50188 21608
rect 50228 21568 50229 21608
rect 50187 21559 50229 21568
rect 50283 21608 50325 21617
rect 50283 21568 50284 21608
rect 50324 21568 50325 21608
rect 50283 21559 50325 21568
rect 50563 21608 50621 21609
rect 50563 21568 50572 21608
rect 50612 21568 50621 21608
rect 50563 21567 50621 21568
rect 50851 21608 50909 21609
rect 50851 21568 50860 21608
rect 50900 21568 50909 21608
rect 50851 21567 50909 21568
rect 50955 21608 50997 21617
rect 50955 21568 50956 21608
rect 50996 21568 50997 21608
rect 50955 21559 50997 21568
rect 51147 21608 51189 21617
rect 51147 21568 51148 21608
rect 51188 21568 51189 21608
rect 51147 21559 51189 21568
rect 52579 21608 52637 21609
rect 52579 21568 52588 21608
rect 52628 21568 52637 21608
rect 52579 21567 52637 21568
rect 52683 21608 52725 21617
rect 52683 21568 52684 21608
rect 52724 21568 52725 21608
rect 52683 21559 52725 21568
rect 3715 21524 3773 21525
rect 2851 21513 2909 21514
rect 2851 21473 2860 21513
rect 2900 21473 2909 21513
rect 3715 21484 3724 21524
rect 3764 21484 3773 21524
rect 3715 21483 3773 21484
rect 5731 21524 5789 21525
rect 5731 21484 5740 21524
rect 5780 21484 5789 21524
rect 5731 21483 5789 21484
rect 5923 21524 5981 21525
rect 5923 21484 5932 21524
rect 5972 21484 5981 21524
rect 5923 21483 5981 21484
rect 26851 21524 26909 21525
rect 26851 21484 26860 21524
rect 26900 21484 26909 21524
rect 26851 21483 26909 21484
rect 27427 21524 27485 21525
rect 27427 21484 27436 21524
rect 27476 21484 27485 21524
rect 27427 21483 27485 21484
rect 48363 21524 48405 21533
rect 48363 21484 48364 21524
rect 48404 21484 48405 21524
rect 48363 21475 48405 21484
rect 2851 21472 2909 21473
rect 5547 21440 5589 21449
rect 5547 21400 5548 21440
rect 5588 21400 5589 21440
rect 5547 21391 5589 21400
rect 26475 21440 26517 21449
rect 26475 21400 26476 21440
rect 26516 21400 26517 21440
rect 26475 21391 26517 21400
rect 27051 21440 27093 21449
rect 27051 21400 27052 21440
rect 27092 21400 27093 21440
rect 27051 21391 27093 21400
rect 27627 21440 27669 21449
rect 27627 21400 27628 21440
rect 27668 21400 27669 21440
rect 27627 21391 27669 21400
rect 29835 21440 29877 21449
rect 29835 21400 29836 21440
rect 29876 21400 29877 21440
rect 29835 21391 29877 21400
rect 32811 21440 32853 21449
rect 32811 21400 32812 21440
rect 32852 21400 32853 21440
rect 32811 21391 32853 21400
rect 33195 21440 33237 21449
rect 33195 21400 33196 21440
rect 33236 21400 33237 21440
rect 33195 21391 33237 21400
rect 35787 21440 35829 21449
rect 35787 21400 35788 21440
rect 35828 21400 35829 21440
rect 35787 21391 35829 21400
rect 36747 21440 36789 21449
rect 36747 21400 36748 21440
rect 36788 21400 36789 21440
rect 36747 21391 36789 21400
rect 39531 21440 39573 21449
rect 39531 21400 39532 21440
rect 39572 21400 39573 21440
rect 39531 21391 39573 21400
rect 49891 21440 49949 21441
rect 49891 21400 49900 21440
rect 49940 21400 49949 21440
rect 49891 21399 49949 21400
rect 51339 21440 51381 21449
rect 51339 21400 51340 21440
rect 51380 21400 51381 21440
rect 51339 21391 51381 21400
rect 2667 21356 2709 21365
rect 2667 21316 2668 21356
rect 2708 21316 2709 21356
rect 2667 21307 2709 21316
rect 3531 21356 3573 21365
rect 3531 21316 3532 21356
rect 3572 21316 3573 21356
rect 3531 21307 3573 21316
rect 6123 21356 6165 21365
rect 6123 21316 6124 21356
rect 6164 21316 6165 21356
rect 6123 21307 6165 21316
rect 28299 21356 28341 21365
rect 28299 21316 28300 21356
rect 28340 21316 28341 21356
rect 28299 21307 28341 21316
rect 28971 21356 29013 21365
rect 28971 21316 28972 21356
rect 29012 21316 29013 21356
rect 28971 21307 29013 21316
rect 45667 21356 45725 21357
rect 45667 21316 45676 21356
rect 45716 21316 45725 21356
rect 45667 21315 45725 21316
rect 48843 21356 48885 21365
rect 48843 21316 48844 21356
rect 48884 21316 48885 21356
rect 48843 21307 48885 21316
rect 576 21188 52800 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 52800 21188
rect 576 21124 52800 21148
rect 31651 21020 31709 21021
rect 31651 20980 31660 21020
rect 31700 20980 31709 21020
rect 31651 20979 31709 20980
rect 46059 21020 46101 21029
rect 46059 20980 46060 21020
rect 46100 20980 46101 21020
rect 46059 20971 46101 20980
rect 46347 21020 46389 21029
rect 46347 20980 46348 21020
rect 46388 20980 46389 21020
rect 46347 20971 46389 20980
rect 50083 21020 50141 21021
rect 50083 20980 50092 21020
rect 50132 20980 50141 21020
rect 50083 20979 50141 20980
rect 52675 21020 52733 21021
rect 52675 20980 52684 21020
rect 52724 20980 52733 21020
rect 52675 20979 52733 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 41739 20936 41781 20945
rect 41739 20896 41740 20936
rect 41780 20896 41781 20936
rect 41739 20887 41781 20896
rect 32035 20852 32093 20853
rect 32035 20812 32044 20852
rect 32084 20812 32093 20852
rect 32035 20811 32093 20812
rect 42883 20852 42941 20853
rect 42883 20812 42892 20852
rect 42932 20812 42941 20852
rect 42883 20811 42941 20812
rect 43459 20852 43517 20853
rect 43459 20812 43468 20852
rect 43508 20812 43517 20852
rect 43459 20811 43517 20812
rect 43651 20852 43709 20853
rect 43651 20812 43660 20852
rect 43700 20812 43709 20852
rect 43651 20811 43709 20812
rect 44131 20852 44189 20853
rect 44131 20812 44140 20852
rect 44180 20812 44189 20852
rect 44131 20811 44189 20812
rect 5443 20768 5501 20769
rect 5443 20728 5452 20768
rect 5492 20728 5501 20768
rect 5443 20727 5501 20728
rect 26947 20768 27005 20769
rect 26947 20728 26956 20768
rect 26996 20728 27005 20768
rect 26947 20727 27005 20728
rect 27811 20768 27869 20769
rect 27811 20728 27820 20768
rect 27860 20728 27869 20768
rect 27811 20727 27869 20728
rect 28203 20768 28245 20777
rect 28203 20728 28204 20768
rect 28244 20728 28245 20768
rect 28203 20719 28245 20728
rect 28683 20768 28725 20777
rect 28683 20728 28684 20768
rect 28724 20728 28725 20768
rect 28683 20719 28725 20728
rect 28875 20768 28917 20777
rect 28875 20728 28876 20768
rect 28916 20728 28917 20768
rect 28875 20719 28917 20728
rect 28963 20768 29021 20769
rect 28963 20728 28972 20768
rect 29012 20728 29021 20768
rect 28963 20727 29021 20728
rect 29635 20768 29693 20769
rect 29635 20728 29644 20768
rect 29684 20728 29693 20768
rect 29635 20727 29693 20728
rect 30499 20768 30557 20769
rect 30499 20728 30508 20768
rect 30548 20728 30557 20768
rect 30499 20727 30557 20728
rect 32707 20768 32765 20769
rect 32707 20728 32716 20768
rect 32756 20728 32765 20768
rect 32707 20727 32765 20728
rect 33571 20768 33629 20769
rect 33571 20728 33580 20768
rect 33620 20728 33629 20768
rect 33571 20727 33629 20728
rect 35779 20768 35837 20769
rect 35779 20728 35788 20768
rect 35828 20728 35837 20768
rect 35779 20727 35837 20728
rect 36643 20768 36701 20769
rect 36643 20728 36652 20768
rect 36692 20728 36701 20768
rect 36643 20727 36701 20728
rect 38275 20768 38333 20769
rect 38275 20728 38284 20768
rect 38324 20728 38333 20768
rect 38275 20727 38333 20728
rect 38379 20768 38421 20777
rect 38379 20728 38380 20768
rect 38420 20728 38421 20768
rect 38379 20719 38421 20728
rect 38571 20768 38613 20777
rect 38571 20728 38572 20768
rect 38612 20728 38613 20768
rect 38571 20719 38613 20728
rect 39139 20768 39197 20769
rect 39139 20728 39148 20768
rect 39188 20728 39197 20768
rect 39139 20727 39197 20728
rect 40003 20768 40061 20769
rect 40003 20728 40012 20768
rect 40052 20728 40061 20768
rect 40003 20727 40061 20728
rect 41923 20768 41981 20769
rect 41923 20728 41932 20768
rect 41972 20728 41981 20768
rect 41923 20727 41981 20728
rect 42027 20768 42069 20777
rect 42027 20728 42028 20768
rect 42068 20728 42069 20768
rect 42027 20719 42069 20728
rect 42219 20768 42261 20777
rect 42219 20728 42220 20768
rect 42260 20728 42261 20768
rect 42219 20719 42261 20728
rect 44811 20768 44853 20777
rect 44811 20728 44812 20768
rect 44852 20728 44853 20768
rect 44811 20719 44853 20728
rect 44907 20768 44949 20777
rect 44907 20728 44908 20768
rect 44948 20728 44949 20768
rect 44907 20719 44949 20728
rect 45003 20768 45045 20777
rect 45003 20728 45004 20768
rect 45044 20728 45045 20768
rect 45003 20719 45045 20728
rect 45099 20768 45141 20777
rect 45099 20728 45100 20768
rect 45140 20728 45141 20768
rect 45099 20719 45141 20728
rect 45483 20768 45525 20777
rect 45483 20728 45484 20768
rect 45524 20728 45525 20768
rect 45483 20719 45525 20728
rect 45675 20768 45717 20777
rect 45675 20728 45676 20768
rect 45716 20728 45717 20768
rect 45675 20719 45717 20728
rect 45763 20768 45821 20769
rect 45763 20728 45772 20768
rect 45812 20728 45821 20768
rect 45763 20727 45821 20728
rect 45963 20768 46005 20777
rect 45963 20728 45964 20768
rect 46004 20728 46005 20768
rect 45963 20719 46005 20728
rect 46147 20768 46205 20769
rect 46147 20728 46156 20768
rect 46196 20728 46205 20768
rect 46147 20727 46205 20728
rect 46347 20768 46389 20777
rect 46347 20728 46348 20768
rect 46388 20728 46389 20768
rect 46347 20719 46389 20728
rect 46539 20768 46581 20777
rect 46539 20728 46540 20768
rect 46580 20728 46581 20768
rect 46539 20719 46581 20728
rect 46627 20768 46685 20769
rect 46627 20728 46636 20768
rect 46676 20728 46685 20768
rect 46627 20727 46685 20728
rect 47691 20768 47733 20777
rect 47691 20728 47692 20768
rect 47732 20728 47733 20768
rect 47691 20719 47733 20728
rect 48067 20768 48125 20769
rect 48067 20728 48076 20768
rect 48116 20728 48125 20768
rect 48067 20727 48125 20728
rect 48931 20768 48989 20769
rect 48931 20728 48940 20768
rect 48980 20728 48989 20768
rect 48931 20727 48989 20728
rect 50283 20768 50325 20777
rect 50283 20728 50284 20768
rect 50324 20728 50325 20768
rect 50283 20719 50325 20728
rect 50659 20768 50717 20769
rect 50659 20728 50668 20768
rect 50708 20728 50717 20768
rect 50659 20727 50717 20728
rect 51523 20768 51581 20769
rect 51523 20728 51532 20768
rect 51572 20728 51581 20768
rect 51523 20727 51581 20728
rect 28779 20684 28821 20693
rect 28779 20644 28780 20684
rect 28820 20644 28821 20684
rect 28779 20635 28821 20644
rect 29259 20684 29301 20693
rect 29259 20644 29260 20684
rect 29300 20644 29301 20684
rect 29259 20635 29301 20644
rect 32331 20684 32373 20693
rect 32331 20644 32332 20684
rect 32372 20644 32373 20684
rect 32331 20635 32373 20644
rect 35403 20684 35445 20693
rect 35403 20644 35404 20684
rect 35444 20644 35445 20684
rect 35403 20635 35445 20644
rect 38763 20684 38805 20693
rect 38763 20644 38764 20684
rect 38804 20644 38805 20684
rect 38763 20635 38805 20644
rect 5547 20600 5589 20609
rect 5547 20560 5548 20600
rect 5588 20560 5589 20600
rect 5547 20551 5589 20560
rect 25795 20600 25853 20601
rect 25795 20560 25804 20600
rect 25844 20560 25853 20600
rect 25795 20559 25853 20560
rect 31851 20600 31893 20609
rect 31851 20560 31852 20600
rect 31892 20560 31893 20600
rect 31851 20551 31893 20560
rect 34723 20600 34781 20601
rect 34723 20560 34732 20600
rect 34772 20560 34781 20600
rect 34723 20559 34781 20560
rect 37795 20600 37853 20601
rect 37795 20560 37804 20600
rect 37844 20560 37853 20600
rect 37795 20559 37853 20560
rect 38467 20600 38525 20601
rect 38467 20560 38476 20600
rect 38516 20560 38525 20600
rect 38467 20559 38525 20560
rect 41155 20600 41213 20601
rect 41155 20560 41164 20600
rect 41204 20560 41213 20600
rect 41155 20559 41213 20560
rect 42115 20600 42173 20601
rect 42115 20560 42124 20600
rect 42164 20560 42173 20600
rect 42115 20559 42173 20560
rect 43083 20600 43125 20609
rect 43083 20560 43084 20600
rect 43124 20560 43125 20600
rect 43083 20551 43125 20560
rect 43275 20600 43317 20609
rect 43275 20560 43276 20600
rect 43316 20560 43317 20600
rect 43275 20551 43317 20560
rect 43851 20600 43893 20609
rect 43851 20560 43852 20600
rect 43892 20560 43893 20600
rect 43851 20551 43893 20560
rect 44331 20600 44373 20609
rect 44331 20560 44332 20600
rect 44372 20560 44373 20600
rect 44331 20551 44373 20560
rect 45571 20600 45629 20601
rect 45571 20560 45580 20600
rect 45620 20560 45629 20600
rect 45571 20559 45629 20560
rect 576 20432 52800 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 52800 20432
rect 576 20368 52800 20392
rect 35683 20264 35741 20265
rect 35683 20224 35692 20264
rect 35732 20224 35741 20264
rect 35683 20223 35741 20224
rect 41163 20180 41205 20189
rect 41163 20140 41164 20180
rect 41204 20140 41205 20180
rect 41163 20131 41205 20140
rect 41451 20180 41493 20189
rect 41451 20140 41452 20180
rect 41492 20140 41493 20180
rect 41451 20131 41493 20140
rect 28982 20109 29024 20118
rect 22731 20096 22773 20105
rect 22731 20056 22732 20096
rect 22772 20056 22773 20096
rect 22731 20047 22773 20056
rect 22827 20096 22869 20105
rect 22827 20056 22828 20096
rect 22868 20056 22869 20096
rect 22827 20047 22869 20056
rect 22923 20096 22965 20105
rect 22923 20056 22924 20096
rect 22964 20056 22965 20096
rect 22923 20047 22965 20056
rect 23019 20096 23061 20105
rect 23019 20056 23020 20096
rect 23060 20056 23061 20096
rect 23019 20047 23061 20056
rect 26667 20096 26709 20105
rect 26667 20056 26668 20096
rect 26708 20056 26709 20096
rect 26667 20047 26709 20056
rect 26859 20096 26901 20105
rect 26859 20056 26860 20096
rect 26900 20056 26901 20096
rect 26859 20047 26901 20056
rect 26947 20096 27005 20097
rect 26947 20056 26956 20096
rect 26996 20056 27005 20096
rect 26947 20055 27005 20056
rect 27907 20096 27965 20097
rect 27907 20056 27916 20096
rect 27956 20056 27965 20096
rect 27907 20055 27965 20056
rect 28203 20096 28245 20105
rect 28203 20056 28204 20096
rect 28244 20056 28245 20096
rect 28203 20047 28245 20056
rect 28299 20096 28341 20105
rect 28299 20056 28300 20096
rect 28340 20056 28341 20096
rect 28299 20047 28341 20056
rect 28779 20096 28821 20105
rect 28779 20056 28780 20096
rect 28820 20056 28821 20096
rect 28779 20047 28821 20056
rect 28875 20096 28917 20105
rect 28875 20056 28876 20096
rect 28916 20056 28917 20096
rect 28982 20069 28983 20109
rect 29023 20069 29024 20109
rect 28982 20060 29024 20069
rect 31171 20096 31229 20097
rect 28875 20047 28917 20056
rect 31171 20056 31180 20096
rect 31220 20056 31229 20096
rect 31171 20055 31229 20056
rect 32043 20096 32085 20105
rect 32043 20056 32044 20096
rect 32084 20056 32085 20096
rect 32043 20047 32085 20056
rect 32619 20096 32661 20105
rect 32619 20056 32620 20096
rect 32660 20056 32661 20096
rect 32619 20047 32661 20056
rect 32715 20096 32757 20105
rect 32715 20056 32716 20096
rect 32756 20056 32757 20096
rect 32715 20047 32757 20056
rect 32811 20096 32853 20105
rect 32811 20056 32812 20096
rect 32852 20056 32853 20096
rect 32811 20047 32853 20056
rect 32907 20096 32949 20105
rect 32907 20056 32908 20096
rect 32948 20056 32949 20096
rect 33283 20096 33341 20097
rect 32907 20047 32949 20056
rect 33099 20081 33141 20090
rect 33099 20041 33100 20081
rect 33140 20041 33141 20081
rect 33283 20056 33292 20096
rect 33332 20056 33341 20096
rect 33283 20055 33341 20056
rect 34915 20096 34973 20097
rect 34915 20056 34924 20096
rect 34964 20056 34973 20096
rect 34915 20055 34973 20056
rect 35019 20096 35061 20105
rect 35019 20056 35020 20096
rect 35060 20056 35061 20096
rect 35019 20047 35061 20056
rect 35211 20096 35253 20105
rect 35211 20056 35212 20096
rect 35252 20056 35253 20096
rect 35211 20047 35253 20056
rect 35491 20096 35549 20097
rect 35491 20056 35500 20096
rect 35540 20056 35549 20096
rect 35491 20055 35549 20056
rect 35595 20096 35637 20105
rect 35595 20056 35596 20096
rect 35636 20056 35637 20096
rect 35595 20047 35637 20056
rect 35787 20096 35829 20105
rect 35787 20056 35788 20096
rect 35828 20056 35829 20096
rect 35787 20047 35829 20056
rect 35979 20096 36021 20105
rect 35979 20056 35980 20096
rect 36020 20056 36021 20096
rect 35979 20047 36021 20056
rect 36075 20096 36117 20105
rect 36075 20056 36076 20096
rect 36116 20056 36117 20096
rect 36075 20047 36117 20056
rect 36171 20096 36213 20105
rect 36171 20056 36172 20096
rect 36212 20056 36213 20096
rect 36171 20047 36213 20056
rect 36267 20096 36309 20105
rect 36267 20056 36268 20096
rect 36308 20056 36309 20096
rect 36267 20047 36309 20056
rect 37515 20096 37557 20105
rect 37515 20056 37516 20096
rect 37556 20056 37557 20096
rect 37515 20047 37557 20056
rect 37699 20096 37757 20097
rect 37699 20056 37708 20096
rect 37748 20056 37757 20096
rect 37699 20055 37757 20056
rect 37891 20096 37949 20097
rect 37891 20056 37900 20096
rect 37940 20056 37949 20096
rect 37891 20055 37949 20056
rect 37995 20096 38037 20105
rect 37995 20056 37996 20096
rect 38036 20056 38037 20096
rect 37995 20047 38037 20056
rect 38187 20096 38229 20105
rect 38187 20056 38188 20096
rect 38228 20056 38229 20096
rect 38187 20047 38229 20056
rect 38563 20096 38621 20097
rect 38563 20056 38572 20096
rect 38612 20056 38621 20096
rect 38563 20055 38621 20056
rect 40963 20096 41021 20097
rect 40963 20056 40972 20096
rect 41012 20056 41021 20096
rect 40963 20055 41021 20056
rect 41067 20096 41109 20105
rect 41067 20056 41068 20096
rect 41108 20056 41109 20096
rect 41067 20047 41109 20056
rect 41259 20096 41301 20105
rect 41259 20056 41260 20096
rect 41300 20056 41301 20096
rect 41259 20047 41301 20056
rect 41827 20096 41885 20097
rect 41827 20056 41836 20096
rect 41876 20056 41885 20096
rect 41827 20055 41885 20056
rect 42691 20096 42749 20097
rect 42691 20056 42700 20096
rect 42740 20056 42749 20096
rect 42691 20055 42749 20056
rect 33099 20032 33141 20041
rect 8995 20012 9053 20013
rect 8995 19972 9004 20012
rect 9044 19972 9053 20012
rect 8995 19971 9053 19972
rect 22339 20012 22397 20013
rect 22339 19972 22348 20012
rect 22388 19972 22397 20012
rect 22339 19971 22397 19972
rect 25603 20012 25661 20013
rect 25603 19972 25612 20012
rect 25652 19972 25661 20012
rect 25603 19971 25661 19972
rect 26275 20012 26333 20013
rect 26275 19972 26284 20012
rect 26324 19972 26333 20012
rect 26275 19971 26333 19972
rect 27139 20012 27197 20013
rect 27139 19972 27148 20012
rect 27188 19972 27197 20012
rect 27139 19971 27197 19972
rect 44323 20012 44381 20013
rect 44323 19972 44332 20012
rect 44372 19972 44381 20012
rect 44323 19971 44381 19972
rect 45283 20012 45341 20013
rect 45283 19972 45292 20012
rect 45332 19972 45341 20012
rect 45283 19971 45341 19972
rect 45667 20012 45725 20013
rect 45667 19972 45676 20012
rect 45716 19972 45725 20012
rect 45667 19971 45725 19972
rect 47491 20012 47549 20013
rect 47491 19972 47500 20012
rect 47540 19972 47549 20012
rect 47491 19971 47549 19972
rect 47875 20012 47933 20013
rect 47875 19972 47884 20012
rect 47924 19972 47933 20012
rect 47875 19971 47933 19972
rect 49315 20012 49373 20013
rect 49315 19972 49324 20012
rect 49364 19972 49373 20012
rect 49315 19971 49373 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 23307 19928 23349 19937
rect 23307 19888 23308 19928
rect 23348 19888 23349 19928
rect 23307 19879 23349 19888
rect 26475 19928 26517 19937
rect 26475 19888 26476 19928
rect 26516 19888 26517 19928
rect 26475 19879 26517 19888
rect 27339 19928 27381 19937
rect 27339 19888 27340 19928
rect 27380 19888 27381 19928
rect 27339 19879 27381 19888
rect 28579 19928 28637 19929
rect 28579 19888 28588 19928
rect 28628 19888 28637 19928
rect 28579 19887 28637 19888
rect 29739 19928 29781 19937
rect 29739 19888 29740 19928
rect 29780 19888 29781 19928
rect 29739 19879 29781 19888
rect 35211 19928 35253 19937
rect 35211 19888 35212 19928
rect 35252 19888 35253 19928
rect 35211 19879 35253 19888
rect 38187 19928 38229 19937
rect 38187 19888 38188 19928
rect 38228 19888 38229 19928
rect 38187 19879 38229 19888
rect 44523 19928 44565 19937
rect 44523 19888 44524 19928
rect 44564 19888 44565 19928
rect 44523 19879 44565 19888
rect 44715 19928 44757 19937
rect 44715 19888 44716 19928
rect 44756 19888 44757 19928
rect 44715 19879 44757 19888
rect 46827 19928 46869 19937
rect 46827 19888 46828 19928
rect 46868 19888 46869 19928
rect 46827 19879 46869 19888
rect 50091 19928 50133 19937
rect 50091 19888 50092 19928
rect 50132 19888 50133 19928
rect 50091 19879 50133 19888
rect 9195 19844 9237 19853
rect 9195 19804 9196 19844
rect 9236 19804 9237 19844
rect 9195 19795 9237 19804
rect 22539 19844 22581 19853
rect 22539 19804 22540 19844
rect 22580 19804 22581 19844
rect 22539 19795 22581 19804
rect 25419 19844 25461 19853
rect 25419 19804 25420 19844
rect 25460 19804 25461 19844
rect 25419 19795 25461 19804
rect 26667 19844 26709 19853
rect 26667 19804 26668 19844
rect 26708 19804 26709 19844
rect 26667 19795 26709 19804
rect 31659 19844 31701 19853
rect 31659 19804 31660 19844
rect 31700 19804 31701 19844
rect 31659 19795 31701 19804
rect 33195 19844 33237 19853
rect 33195 19804 33196 19844
rect 33236 19804 33237 19844
rect 33195 19795 33237 19804
rect 37611 19844 37653 19853
rect 37611 19804 37612 19844
rect 37652 19804 37653 19844
rect 37611 19795 37653 19804
rect 40107 19844 40149 19853
rect 40107 19804 40108 19844
rect 40148 19804 40149 19844
rect 40107 19795 40149 19804
rect 43843 19844 43901 19845
rect 43843 19804 43852 19844
rect 43892 19804 43901 19844
rect 43843 19803 43901 19804
rect 45099 19844 45141 19853
rect 45099 19804 45100 19844
rect 45140 19804 45141 19844
rect 45099 19795 45141 19804
rect 45483 19844 45525 19853
rect 45483 19804 45484 19844
rect 45524 19804 45525 19844
rect 45483 19795 45525 19804
rect 47307 19844 47349 19853
rect 47307 19804 47308 19844
rect 47348 19804 47349 19844
rect 47307 19795 47349 19804
rect 47691 19844 47733 19853
rect 47691 19804 47692 19844
rect 47732 19804 47733 19844
rect 47691 19795 47733 19804
rect 49131 19844 49173 19853
rect 49131 19804 49132 19844
rect 49172 19804 49173 19844
rect 49131 19795 49173 19804
rect 576 19676 52800 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 52800 19676
rect 576 19612 52800 19636
rect 11683 19508 11741 19509
rect 11683 19468 11692 19508
rect 11732 19468 11741 19508
rect 11683 19467 11741 19468
rect 22155 19508 22197 19517
rect 22155 19468 22156 19508
rect 22196 19468 22197 19508
rect 22155 19459 22197 19468
rect 32427 19508 32469 19517
rect 32427 19468 32428 19508
rect 32468 19468 32469 19508
rect 32427 19459 32469 19468
rect 32899 19508 32957 19509
rect 32899 19468 32908 19508
rect 32948 19468 32957 19508
rect 32899 19467 32957 19468
rect 35787 19508 35829 19517
rect 35787 19468 35788 19508
rect 35828 19468 35829 19508
rect 35787 19459 35829 19468
rect 39043 19508 39101 19509
rect 39043 19468 39052 19508
rect 39092 19468 39101 19508
rect 39043 19467 39101 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 6603 19424 6645 19433
rect 6603 19384 6604 19424
rect 6644 19384 6645 19424
rect 6603 19375 6645 19384
rect 8811 19424 8853 19433
rect 8811 19384 8812 19424
rect 8852 19384 8853 19424
rect 8811 19375 8853 19384
rect 25899 19424 25941 19433
rect 25899 19384 25900 19424
rect 25940 19384 25941 19424
rect 25899 19375 25941 19384
rect 33867 19424 33909 19433
rect 33867 19384 33868 19424
rect 33908 19384 33909 19424
rect 33867 19375 33909 19384
rect 36067 19424 36125 19425
rect 36067 19384 36076 19424
rect 36116 19384 36125 19424
rect 36067 19383 36125 19384
rect 38283 19424 38325 19433
rect 38283 19384 38284 19424
rect 38324 19384 38325 19424
rect 38283 19375 38325 19384
rect 40299 19424 40341 19433
rect 40299 19384 40300 19424
rect 40340 19384 40341 19424
rect 40299 19375 40341 19384
rect 40683 19424 40725 19433
rect 40683 19384 40684 19424
rect 40724 19384 40725 19424
rect 40683 19375 40725 19384
rect 43555 19424 43613 19425
rect 43555 19384 43564 19424
rect 43604 19384 43613 19424
rect 43555 19383 43613 19384
rect 21571 19340 21629 19341
rect 21571 19300 21580 19340
rect 21620 19300 21629 19340
rect 21571 19299 21629 19300
rect 21955 19340 22013 19341
rect 21955 19300 21964 19340
rect 22004 19300 22013 19340
rect 21955 19299 22013 19300
rect 37219 19340 37277 19341
rect 37219 19300 37228 19340
rect 37268 19300 37277 19340
rect 37219 19299 37277 19300
rect 41251 19340 41309 19341
rect 41251 19300 41260 19340
rect 41300 19300 41309 19340
rect 41251 19299 41309 19300
rect 41635 19340 41693 19341
rect 41635 19300 41644 19340
rect 41684 19300 41693 19340
rect 41635 19299 41693 19300
rect 42019 19340 42077 19341
rect 42019 19300 42028 19340
rect 42068 19300 42077 19340
rect 42019 19299 42077 19300
rect 8331 19256 8373 19265
rect 8331 19216 8332 19256
rect 8372 19216 8373 19256
rect 8331 19207 8373 19216
rect 8523 19256 8565 19265
rect 8523 19216 8524 19256
rect 8564 19216 8565 19256
rect 8523 19207 8565 19216
rect 8611 19256 8669 19257
rect 8611 19216 8620 19256
rect 8660 19216 8669 19256
rect 8611 19215 8669 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 9003 19256 9045 19265
rect 9003 19216 9004 19256
rect 9044 19216 9045 19256
rect 9003 19207 9045 19216
rect 9091 19256 9149 19257
rect 9091 19216 9100 19256
rect 9140 19216 9149 19256
rect 9091 19215 9149 19216
rect 9291 19256 9333 19265
rect 9291 19216 9292 19256
rect 9332 19216 9333 19256
rect 9291 19207 9333 19216
rect 9667 19256 9725 19257
rect 9667 19216 9676 19256
rect 9716 19216 9725 19256
rect 9667 19215 9725 19216
rect 10531 19256 10589 19257
rect 10531 19216 10540 19256
rect 10580 19216 10589 19256
rect 10531 19215 10589 19216
rect 22339 19256 22397 19257
rect 22339 19216 22348 19256
rect 22388 19216 22397 19256
rect 22339 19215 22397 19216
rect 22443 19256 22485 19265
rect 22443 19216 22444 19256
rect 22484 19216 22485 19256
rect 23203 19256 23261 19257
rect 22443 19207 22485 19216
rect 22635 19242 22677 19251
rect 22635 19202 22636 19242
rect 22676 19202 22677 19242
rect 23203 19216 23212 19256
rect 23252 19216 23261 19256
rect 23203 19215 23261 19216
rect 24067 19256 24125 19257
rect 24067 19216 24076 19256
rect 24116 19216 24125 19256
rect 24067 19215 24125 19216
rect 26467 19256 26525 19257
rect 26467 19216 26476 19256
rect 26516 19216 26525 19256
rect 26467 19215 26525 19216
rect 27372 19256 27414 19265
rect 27372 19216 27373 19256
rect 27413 19216 27414 19256
rect 27372 19207 27414 19216
rect 29635 19256 29693 19257
rect 29635 19216 29644 19256
rect 29684 19216 29693 19256
rect 29635 19215 29693 19216
rect 30499 19256 30557 19257
rect 30499 19216 30508 19256
rect 30548 19216 30557 19256
rect 30499 19215 30557 19216
rect 32131 19256 32189 19257
rect 32131 19216 32140 19256
rect 32180 19216 32189 19256
rect 32131 19215 32189 19216
rect 32235 19256 32277 19265
rect 32235 19216 32236 19256
rect 32276 19216 32277 19256
rect 32235 19207 32277 19216
rect 32427 19256 32469 19265
rect 32427 19216 32428 19256
rect 32468 19216 32469 19256
rect 32427 19207 32469 19216
rect 33195 19256 33237 19265
rect 33195 19216 33196 19256
rect 33236 19216 33237 19256
rect 33195 19207 33237 19216
rect 33291 19256 33333 19265
rect 33291 19216 33292 19256
rect 33332 19216 33333 19256
rect 33291 19207 33333 19216
rect 33571 19256 33629 19257
rect 33571 19216 33580 19256
rect 33620 19216 33629 19256
rect 33571 19215 33629 19216
rect 35683 19256 35741 19257
rect 35683 19216 35692 19256
rect 35732 19216 35741 19256
rect 35683 19215 35741 19216
rect 35883 19256 35925 19265
rect 35883 19216 35884 19256
rect 35924 19216 35925 19256
rect 35883 19207 35925 19216
rect 36363 19256 36405 19265
rect 36363 19216 36364 19256
rect 36404 19216 36405 19256
rect 36363 19207 36405 19216
rect 36459 19256 36501 19265
rect 36459 19216 36460 19256
rect 36500 19216 36501 19256
rect 36459 19207 36501 19216
rect 36739 19256 36797 19257
rect 36739 19216 36748 19256
rect 36788 19216 36797 19256
rect 36739 19215 36797 19216
rect 38179 19256 38237 19257
rect 38179 19216 38188 19256
rect 38228 19216 38237 19256
rect 38179 19215 38237 19216
rect 38379 19256 38421 19265
rect 38379 19216 38380 19256
rect 38420 19216 38421 19256
rect 38379 19207 38421 19216
rect 38563 19256 38621 19257
rect 38563 19216 38572 19256
rect 38612 19216 38621 19256
rect 38563 19215 38621 19216
rect 38667 19256 38709 19265
rect 38667 19216 38668 19256
rect 38708 19216 38709 19256
rect 38667 19207 38709 19216
rect 38859 19256 38901 19265
rect 38859 19216 38860 19256
rect 38900 19216 38901 19256
rect 38859 19207 38901 19216
rect 39339 19256 39381 19265
rect 39339 19216 39340 19256
rect 39380 19216 39381 19256
rect 39339 19207 39381 19216
rect 39435 19256 39477 19265
rect 39435 19216 39436 19256
rect 39476 19216 39477 19256
rect 39435 19207 39477 19216
rect 39715 19256 39773 19257
rect 39715 19216 39724 19256
rect 39764 19216 39773 19256
rect 39715 19215 39773 19216
rect 42219 19256 42261 19265
rect 42219 19216 42220 19256
rect 42260 19216 42261 19256
rect 42219 19207 42261 19216
rect 42315 19256 42357 19265
rect 42315 19216 42316 19256
rect 42356 19216 42357 19256
rect 42315 19207 42357 19216
rect 42411 19256 42453 19265
rect 42411 19216 42412 19256
rect 42452 19216 42453 19256
rect 42411 19207 42453 19216
rect 42507 19256 42549 19265
rect 42507 19216 42508 19256
rect 42548 19216 42549 19256
rect 42507 19207 42549 19216
rect 42883 19256 42941 19257
rect 42883 19216 42892 19256
rect 42932 19216 42941 19256
rect 43275 19256 43317 19265
rect 42883 19215 42941 19216
rect 43179 19229 43221 19238
rect 22635 19193 22677 19202
rect 43179 19189 43180 19229
rect 43220 19189 43221 19229
rect 43275 19216 43276 19256
rect 43316 19216 43317 19256
rect 43275 19207 43317 19216
rect 44131 19256 44189 19257
rect 44131 19216 44140 19256
rect 44180 19216 44189 19256
rect 44131 19215 44189 19216
rect 44995 19256 45053 19257
rect 44995 19216 45004 19256
rect 45044 19216 45053 19256
rect 44995 19215 45053 19216
rect 46723 19256 46781 19257
rect 46723 19216 46732 19256
rect 46772 19216 46781 19256
rect 46723 19215 46781 19216
rect 47587 19256 47645 19257
rect 47587 19216 47596 19256
rect 47636 19216 47645 19256
rect 47587 19215 47645 19216
rect 49035 19256 49077 19265
rect 49035 19216 49036 19256
rect 49076 19216 49077 19256
rect 49035 19207 49077 19216
rect 49227 19256 49269 19265
rect 49227 19216 49228 19256
rect 49268 19216 49269 19256
rect 49227 19207 49269 19216
rect 49315 19256 49373 19257
rect 49315 19216 49324 19256
rect 49364 19216 49373 19256
rect 49315 19215 49373 19216
rect 49987 19256 50045 19257
rect 49987 19216 49996 19256
rect 50036 19216 50045 19256
rect 49987 19215 50045 19216
rect 50851 19256 50909 19257
rect 50851 19216 50860 19256
rect 50900 19216 50909 19256
rect 50851 19215 50909 19216
rect 22827 19172 22869 19181
rect 22827 19132 22828 19172
rect 22868 19132 22869 19172
rect 22827 19123 22869 19132
rect 26091 19172 26133 19181
rect 26091 19132 26092 19172
rect 26132 19132 26133 19172
rect 26091 19123 26133 19132
rect 29259 19172 29301 19181
rect 43179 19180 43221 19189
rect 29259 19132 29260 19172
rect 29300 19132 29301 19172
rect 29259 19123 29301 19132
rect 43755 19172 43797 19181
rect 43755 19132 43756 19172
rect 43796 19132 43797 19172
rect 43755 19123 43797 19132
rect 46347 19172 46389 19181
rect 46347 19132 46348 19172
rect 46388 19132 46389 19172
rect 46347 19123 46389 19132
rect 49131 19172 49173 19181
rect 49131 19132 49132 19172
rect 49172 19132 49173 19172
rect 49131 19123 49173 19132
rect 49611 19172 49653 19181
rect 49611 19132 49612 19172
rect 49652 19132 49653 19172
rect 49611 19123 49653 19132
rect 8419 19088 8477 19089
rect 8419 19048 8428 19088
rect 8468 19048 8477 19088
rect 8419 19047 8477 19048
rect 11683 19088 11741 19089
rect 11683 19048 11692 19088
rect 11732 19048 11741 19088
rect 11683 19047 11741 19048
rect 21771 19088 21813 19097
rect 21771 19048 21772 19088
rect 21812 19048 21813 19088
rect 21771 19039 21813 19048
rect 22155 19088 22197 19097
rect 22155 19048 22156 19088
rect 22196 19048 22197 19088
rect 22155 19039 22197 19048
rect 22531 19088 22589 19089
rect 22531 19048 22540 19088
rect 22580 19048 22589 19088
rect 22531 19047 22589 19048
rect 25219 19088 25277 19089
rect 25219 19048 25228 19088
rect 25268 19048 25277 19088
rect 25219 19047 25277 19048
rect 28483 19088 28541 19089
rect 28483 19048 28492 19088
rect 28532 19048 28541 19088
rect 28483 19047 28541 19048
rect 31651 19088 31709 19089
rect 31651 19048 31660 19088
rect 31700 19048 31709 19088
rect 31651 19047 31709 19048
rect 37035 19088 37077 19097
rect 37035 19048 37036 19088
rect 37076 19048 37077 19088
rect 37035 19039 37077 19048
rect 38755 19088 38813 19089
rect 38755 19048 38764 19088
rect 38804 19048 38813 19088
rect 38755 19047 38813 19048
rect 41067 19088 41109 19097
rect 41067 19048 41068 19088
rect 41108 19048 41109 19088
rect 41067 19039 41109 19048
rect 41451 19088 41493 19097
rect 41451 19048 41452 19088
rect 41492 19048 41493 19088
rect 41451 19039 41493 19048
rect 41835 19088 41877 19097
rect 41835 19048 41836 19088
rect 41876 19048 41877 19088
rect 41835 19039 41877 19048
rect 46147 19088 46205 19089
rect 46147 19048 46156 19088
rect 46196 19048 46205 19088
rect 46147 19047 46205 19048
rect 48739 19088 48797 19089
rect 48739 19048 48748 19088
rect 48788 19048 48797 19088
rect 48739 19047 48797 19048
rect 52003 19088 52061 19089
rect 52003 19048 52012 19088
rect 52052 19048 52061 19088
rect 52003 19047 52061 19048
rect 576 18920 52800 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 52800 18920
rect 576 18856 52800 18880
rect 9003 18752 9045 18761
rect 9003 18712 9004 18752
rect 9044 18712 9045 18752
rect 9003 18703 9045 18712
rect 26083 18752 26141 18753
rect 26083 18712 26092 18752
rect 26132 18712 26141 18752
rect 26083 18711 26141 18712
rect 29347 18752 29405 18753
rect 29347 18712 29356 18752
rect 29396 18712 29405 18752
rect 29347 18711 29405 18712
rect 42891 18752 42933 18761
rect 42891 18712 42892 18752
rect 42932 18712 42933 18752
rect 42891 18703 42933 18712
rect 44035 18752 44093 18753
rect 44035 18712 44044 18752
rect 44084 18712 44093 18752
rect 44035 18711 44093 18712
rect 8331 18668 8373 18677
rect 8331 18628 8332 18668
rect 8372 18628 8373 18668
rect 8331 18619 8373 18628
rect 8811 18668 8853 18677
rect 8811 18628 8812 18668
rect 8852 18628 8853 18668
rect 8811 18619 8853 18628
rect 9483 18668 9525 18677
rect 9483 18628 9484 18668
rect 9524 18628 9525 18668
rect 9483 18619 9525 18628
rect 23115 18668 23157 18677
rect 23115 18628 23116 18668
rect 23156 18628 23157 18668
rect 23115 18619 23157 18628
rect 30603 18668 30645 18677
rect 30603 18628 30604 18668
rect 30644 18628 30645 18668
rect 30603 18619 30645 18628
rect 32619 18668 32661 18677
rect 32619 18628 32620 18668
rect 32660 18628 32661 18668
rect 32619 18619 32661 18628
rect 35787 18668 35829 18677
rect 35787 18628 35788 18668
rect 35828 18628 35829 18668
rect 35787 18619 35829 18628
rect 36171 18668 36213 18677
rect 36171 18628 36172 18668
rect 36212 18628 36213 18668
rect 36171 18619 36213 18628
rect 38763 18668 38805 18677
rect 38763 18628 38764 18668
rect 38804 18628 38805 18668
rect 38763 18619 38805 18628
rect 48075 18668 48117 18677
rect 48075 18628 48076 18668
rect 48116 18628 48117 18668
rect 48075 18619 48117 18628
rect 48651 18668 48693 18677
rect 48651 18628 48652 18668
rect 48692 18628 48693 18668
rect 48651 18619 48693 18628
rect 49419 18668 49461 18677
rect 49419 18628 49420 18668
rect 49460 18628 49461 18668
rect 49419 18619 49461 18628
rect 7075 18584 7133 18585
rect 7075 18544 7084 18584
rect 7124 18544 7133 18584
rect 7075 18543 7133 18544
rect 7939 18584 7997 18585
rect 7939 18544 7948 18584
rect 7988 18544 7997 18584
rect 7939 18543 7997 18544
rect 8523 18584 8565 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8523 18535 8565 18544
rect 8715 18584 8757 18593
rect 8715 18544 8716 18584
rect 8756 18544 8757 18584
rect 8611 18542 8669 18543
rect 8611 18502 8620 18542
rect 8660 18502 8669 18542
rect 8715 18535 8757 18544
rect 9379 18584 9437 18585
rect 9379 18544 9388 18584
rect 9428 18544 9437 18584
rect 9379 18543 9437 18544
rect 9579 18584 9621 18593
rect 9579 18544 9580 18584
rect 9620 18544 9621 18584
rect 9579 18535 9621 18544
rect 22723 18584 22781 18585
rect 22723 18544 22732 18584
rect 22772 18544 22781 18584
rect 22723 18543 22781 18544
rect 23019 18584 23061 18593
rect 23019 18544 23020 18584
rect 23060 18544 23061 18584
rect 23019 18535 23061 18544
rect 25315 18584 25373 18585
rect 25315 18544 25324 18584
rect 25364 18544 25373 18584
rect 25315 18543 25373 18544
rect 25419 18584 25461 18593
rect 25419 18544 25420 18584
rect 25460 18544 25461 18584
rect 25419 18535 25461 18544
rect 25611 18584 25653 18593
rect 25611 18544 25612 18584
rect 25652 18544 25653 18584
rect 25611 18535 25653 18544
rect 25891 18584 25949 18585
rect 25891 18544 25900 18584
rect 25940 18544 25949 18584
rect 25891 18543 25949 18544
rect 25995 18584 26037 18593
rect 25995 18544 25996 18584
rect 26036 18544 26037 18584
rect 25995 18535 26037 18544
rect 26187 18584 26229 18593
rect 26187 18544 26188 18584
rect 26228 18544 26229 18584
rect 26187 18535 26229 18544
rect 26379 18584 26421 18593
rect 26379 18544 26380 18584
rect 26420 18544 26421 18584
rect 26379 18535 26421 18544
rect 26475 18584 26517 18593
rect 26475 18544 26476 18584
rect 26516 18544 26517 18584
rect 26475 18535 26517 18544
rect 26571 18584 26613 18593
rect 26571 18544 26572 18584
rect 26612 18544 26613 18584
rect 26571 18535 26613 18544
rect 26667 18584 26709 18593
rect 26667 18544 26668 18584
rect 26708 18544 26709 18584
rect 26667 18535 26709 18544
rect 28675 18584 28733 18585
rect 28675 18544 28684 18584
rect 28724 18544 28733 18584
rect 28675 18543 28733 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 28779 18535 28821 18544
rect 28971 18584 29013 18593
rect 28971 18544 28972 18584
rect 29012 18544 29013 18584
rect 28971 18535 29013 18544
rect 29155 18584 29213 18585
rect 29155 18544 29164 18584
rect 29204 18544 29213 18584
rect 29155 18543 29213 18544
rect 29259 18584 29301 18593
rect 29259 18544 29260 18584
rect 29300 18544 29301 18584
rect 29259 18535 29301 18544
rect 29451 18584 29493 18593
rect 29451 18544 29452 18584
rect 29492 18544 29493 18584
rect 29451 18535 29493 18544
rect 29643 18584 29685 18593
rect 29643 18544 29644 18584
rect 29684 18544 29685 18584
rect 29643 18535 29685 18544
rect 29739 18584 29781 18593
rect 29739 18544 29740 18584
rect 29780 18544 29781 18584
rect 29739 18535 29781 18544
rect 29835 18584 29877 18593
rect 29835 18544 29836 18584
rect 29876 18544 29877 18584
rect 29835 18535 29877 18544
rect 29931 18584 29973 18593
rect 29931 18544 29932 18584
rect 29972 18544 29973 18584
rect 29931 18535 29973 18544
rect 30211 18584 30269 18585
rect 30211 18544 30220 18584
rect 30260 18544 30269 18584
rect 30211 18543 30269 18544
rect 30507 18584 30549 18593
rect 30507 18544 30508 18584
rect 30548 18544 30549 18584
rect 30507 18535 30549 18544
rect 31083 18584 31125 18593
rect 31083 18544 31084 18584
rect 31124 18544 31125 18584
rect 31083 18535 31125 18544
rect 31267 18584 31325 18585
rect 31267 18544 31276 18584
rect 31316 18544 31325 18584
rect 31267 18543 31325 18544
rect 31843 18584 31901 18585
rect 31843 18544 31852 18584
rect 31892 18544 31901 18584
rect 31843 18543 31901 18544
rect 31947 18584 31989 18593
rect 31947 18544 31948 18584
rect 31988 18544 31989 18584
rect 31947 18535 31989 18544
rect 32139 18584 32181 18593
rect 32139 18544 32140 18584
rect 32180 18544 32181 18584
rect 32139 18535 32181 18544
rect 32523 18584 32565 18593
rect 32523 18544 32524 18584
rect 32564 18544 32565 18584
rect 32523 18535 32565 18544
rect 32715 18584 32757 18593
rect 32715 18544 32716 18584
rect 32756 18544 32757 18584
rect 32715 18535 32757 18544
rect 32803 18584 32861 18585
rect 32803 18544 32812 18584
rect 32852 18544 32861 18584
rect 32803 18543 32861 18544
rect 33003 18584 33045 18593
rect 33003 18544 33004 18584
rect 33044 18544 33045 18584
rect 33003 18535 33045 18544
rect 33379 18584 33437 18585
rect 33379 18544 33388 18584
rect 33428 18544 33437 18584
rect 33379 18543 33437 18544
rect 34243 18584 34301 18585
rect 34243 18544 34252 18584
rect 34292 18544 34301 18584
rect 34243 18543 34301 18544
rect 35691 18584 35733 18593
rect 35691 18544 35692 18584
rect 35732 18544 35733 18584
rect 35691 18535 35733 18544
rect 35883 18584 35925 18593
rect 35883 18544 35884 18584
rect 35924 18544 35925 18584
rect 35883 18535 35925 18544
rect 35971 18584 36029 18585
rect 35971 18544 35980 18584
rect 36020 18544 36029 18584
rect 35971 18543 36029 18544
rect 36547 18584 36605 18585
rect 36547 18544 36556 18584
rect 36596 18544 36605 18584
rect 36547 18543 36605 18544
rect 37411 18584 37469 18585
rect 37411 18544 37420 18584
rect 37460 18544 37469 18584
rect 37411 18543 37469 18544
rect 39139 18584 39197 18585
rect 39139 18544 39148 18584
rect 39188 18544 39197 18584
rect 39139 18543 39197 18544
rect 39963 18584 40005 18593
rect 39963 18544 39964 18584
rect 40004 18544 40005 18584
rect 39963 18535 40005 18544
rect 41931 18584 41973 18593
rect 41931 18544 41932 18584
rect 41972 18544 41973 18584
rect 41931 18535 41973 18544
rect 42123 18584 42165 18593
rect 42123 18544 42124 18584
rect 42164 18544 42165 18584
rect 42123 18535 42165 18544
rect 42211 18584 42269 18585
rect 42211 18544 42220 18584
rect 42260 18544 42269 18584
rect 42211 18543 42269 18544
rect 42411 18584 42453 18593
rect 42411 18544 42412 18584
rect 42452 18544 42453 18584
rect 42411 18535 42453 18544
rect 42603 18584 42645 18593
rect 42603 18544 42604 18584
rect 42644 18544 42645 18584
rect 42603 18535 42645 18544
rect 42691 18584 42749 18585
rect 42691 18544 42700 18584
rect 42740 18544 42749 18584
rect 42691 18543 42749 18544
rect 43563 18584 43605 18593
rect 43563 18544 43564 18584
rect 43604 18544 43605 18584
rect 43563 18535 43605 18544
rect 43659 18584 43701 18593
rect 43659 18544 43660 18584
rect 43700 18544 43701 18584
rect 43659 18535 43701 18544
rect 43747 18584 43805 18585
rect 43747 18544 43756 18584
rect 43796 18544 43805 18584
rect 43747 18543 43805 18544
rect 43947 18584 43989 18593
rect 43947 18544 43948 18584
rect 43988 18544 43989 18584
rect 43947 18535 43989 18544
rect 44139 18584 44181 18593
rect 44139 18544 44140 18584
rect 44180 18544 44181 18584
rect 44139 18535 44181 18544
rect 44227 18584 44285 18585
rect 44227 18544 44236 18584
rect 44276 18544 44285 18584
rect 44227 18543 44285 18544
rect 44419 18584 44477 18585
rect 44419 18544 44428 18584
rect 44468 18544 44477 18584
rect 44419 18543 44477 18544
rect 44523 18584 44565 18593
rect 44523 18544 44524 18584
rect 44564 18544 44565 18584
rect 44523 18535 44565 18544
rect 44619 18584 44661 18593
rect 44619 18544 44620 18584
rect 44660 18544 44661 18584
rect 44619 18535 44661 18544
rect 46155 18584 46197 18593
rect 46155 18544 46156 18584
rect 46196 18544 46197 18584
rect 46155 18535 46197 18544
rect 46339 18584 46397 18585
rect 46339 18544 46348 18584
rect 46388 18544 46397 18584
rect 46339 18543 46397 18544
rect 46723 18584 46781 18585
rect 46723 18544 46732 18584
rect 46772 18544 46781 18584
rect 46723 18543 46781 18544
rect 46827 18584 46869 18593
rect 46827 18544 46828 18584
rect 46868 18544 46869 18584
rect 46827 18535 46869 18544
rect 47019 18584 47061 18593
rect 47019 18544 47020 18584
rect 47060 18544 47061 18584
rect 47019 18535 47061 18544
rect 47403 18584 47445 18593
rect 47403 18544 47404 18584
rect 47444 18544 47445 18584
rect 47403 18535 47445 18544
rect 47499 18584 47541 18593
rect 47499 18544 47500 18584
rect 47540 18544 47541 18584
rect 47499 18535 47541 18544
rect 47595 18584 47637 18593
rect 47595 18544 47596 18584
rect 47636 18544 47637 18584
rect 47595 18535 47637 18544
rect 47691 18584 47733 18593
rect 47691 18544 47692 18584
rect 47732 18544 47733 18584
rect 47691 18535 47733 18544
rect 47971 18584 48029 18585
rect 47971 18544 47980 18584
rect 48020 18544 48029 18584
rect 47971 18543 48029 18544
rect 48171 18584 48213 18593
rect 48171 18544 48172 18584
rect 48212 18544 48213 18584
rect 48171 18535 48213 18544
rect 48747 18584 48789 18593
rect 48747 18544 48748 18584
rect 48788 18544 48789 18584
rect 48747 18535 48789 18544
rect 49027 18584 49085 18585
rect 49027 18544 49036 18584
rect 49076 18544 49085 18584
rect 49027 18543 49085 18544
rect 49315 18584 49373 18585
rect 49315 18544 49324 18584
rect 49364 18544 49373 18584
rect 49315 18543 49373 18544
rect 49515 18584 49557 18593
rect 49515 18544 49516 18584
rect 49556 18544 49557 18584
rect 49515 18535 49557 18544
rect 52291 18584 52349 18585
rect 52291 18544 52300 18584
rect 52340 18544 52349 18584
rect 52291 18543 52349 18544
rect 52675 18584 52733 18585
rect 52675 18544 52684 18584
rect 52724 18544 52733 18584
rect 52675 18543 52733 18544
rect 8611 18501 8669 18502
rect 9187 18500 9245 18501
rect 9187 18460 9196 18500
rect 9236 18460 9245 18500
rect 9187 18459 9245 18460
rect 21475 18500 21533 18501
rect 21475 18460 21484 18500
rect 21524 18460 21533 18500
rect 21475 18459 21533 18460
rect 22051 18500 22109 18501
rect 22051 18460 22060 18500
rect 22100 18460 22109 18500
rect 22051 18459 22109 18460
rect 22243 18500 22301 18501
rect 22243 18460 22252 18500
rect 22292 18460 22301 18500
rect 22243 18459 22301 18460
rect 23587 18500 23645 18501
rect 23587 18460 23596 18500
rect 23636 18460 23645 18500
rect 23587 18459 23645 18460
rect 23971 18500 24029 18501
rect 23971 18460 23980 18500
rect 24020 18460 24029 18500
rect 23971 18459 24029 18460
rect 24355 18500 24413 18501
rect 24355 18460 24364 18500
rect 24404 18460 24413 18500
rect 24355 18459 24413 18460
rect 41163 18500 41205 18509
rect 41163 18460 41164 18500
rect 41204 18460 41205 18500
rect 41163 18451 41205 18460
rect 41731 18500 41789 18501
rect 41731 18460 41740 18500
rect 41780 18460 41789 18500
rect 41731 18459 41789 18460
rect 43075 18500 43133 18501
rect 43075 18460 43084 18500
rect 43124 18460 43133 18500
rect 43075 18459 43133 18460
rect 49891 18500 49949 18501
rect 49891 18460 49900 18500
rect 49940 18460 49949 18500
rect 49891 18459 49949 18460
rect 50563 18500 50621 18501
rect 50563 18460 50572 18500
rect 50612 18460 50621 18500
rect 50563 18459 50621 18460
rect 51331 18500 51389 18501
rect 51331 18460 51340 18500
rect 51380 18460 51389 18500
rect 51331 18459 51389 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 9771 18416 9813 18425
rect 9771 18376 9772 18416
rect 9812 18376 9813 18416
rect 9771 18367 9813 18376
rect 23787 18416 23829 18425
rect 23787 18376 23788 18416
rect 23828 18376 23829 18416
rect 23787 18367 23829 18376
rect 25611 18416 25653 18425
rect 25611 18376 25612 18416
rect 25652 18376 25653 18416
rect 25611 18367 25653 18376
rect 28971 18416 29013 18425
rect 28971 18376 28972 18416
rect 29012 18376 29013 18416
rect 28971 18367 29013 18376
rect 30883 18416 30941 18417
rect 30883 18376 30892 18416
rect 30932 18376 30941 18416
rect 30883 18375 30941 18376
rect 32139 18416 32181 18425
rect 32139 18376 32140 18416
rect 32180 18376 32181 18416
rect 32139 18367 32181 18376
rect 42411 18416 42453 18425
rect 42411 18376 42412 18416
rect 42452 18376 42453 18416
rect 42411 18367 42453 18376
rect 46251 18416 46293 18425
rect 46251 18376 46252 18416
rect 46292 18376 46293 18416
rect 46251 18367 46293 18376
rect 48355 18416 48413 18417
rect 48355 18376 48364 18416
rect 48404 18376 48413 18416
rect 48355 18375 48413 18376
rect 50763 18416 50805 18425
rect 50763 18376 50764 18416
rect 50804 18376 50805 18416
rect 50763 18367 50805 18376
rect 5923 18332 5981 18333
rect 5923 18292 5932 18332
rect 5972 18292 5981 18332
rect 5923 18291 5981 18292
rect 9003 18332 9045 18341
rect 9003 18292 9004 18332
rect 9044 18292 9045 18332
rect 9003 18283 9045 18292
rect 21675 18332 21717 18341
rect 21675 18292 21676 18332
rect 21716 18292 21717 18332
rect 21675 18283 21717 18292
rect 21867 18332 21909 18341
rect 21867 18292 21868 18332
rect 21908 18292 21909 18332
rect 21867 18283 21909 18292
rect 22443 18332 22485 18341
rect 22443 18292 22444 18332
rect 22484 18292 22485 18332
rect 22443 18283 22485 18292
rect 23395 18332 23453 18333
rect 23395 18292 23404 18332
rect 23444 18292 23453 18332
rect 23395 18291 23453 18292
rect 24171 18332 24213 18341
rect 24171 18292 24172 18332
rect 24212 18292 24213 18332
rect 24171 18283 24213 18292
rect 24555 18332 24597 18341
rect 24555 18292 24556 18332
rect 24596 18292 24597 18332
rect 24555 18283 24597 18292
rect 31179 18332 31221 18341
rect 31179 18292 31180 18332
rect 31220 18292 31221 18332
rect 31179 18283 31221 18292
rect 35395 18332 35453 18333
rect 35395 18292 35404 18332
rect 35444 18292 35453 18332
rect 35395 18291 35453 18292
rect 38563 18332 38621 18333
rect 38563 18292 38572 18332
rect 38612 18292 38621 18332
rect 38563 18291 38621 18292
rect 41547 18332 41589 18341
rect 41547 18292 41548 18332
rect 41588 18292 41589 18332
rect 41547 18283 41589 18292
rect 41931 18332 41973 18341
rect 41931 18292 41932 18332
rect 41972 18292 41973 18332
rect 41931 18283 41973 18292
rect 42891 18332 42933 18341
rect 42891 18292 42892 18332
rect 42932 18292 42933 18332
rect 42891 18283 42933 18292
rect 47019 18332 47061 18341
rect 47019 18292 47020 18332
rect 47060 18292 47061 18332
rect 47019 18283 47061 18292
rect 50091 18332 50133 18341
rect 50091 18292 50092 18332
rect 50132 18292 50133 18332
rect 50091 18283 50133 18292
rect 50379 18332 50421 18341
rect 50379 18292 50380 18332
rect 50420 18292 50421 18332
rect 50379 18283 50421 18292
rect 51147 18332 51189 18341
rect 51147 18292 51148 18332
rect 51188 18292 51189 18332
rect 51147 18283 51189 18292
rect 52395 18332 52437 18341
rect 52395 18292 52396 18332
rect 52436 18292 52437 18332
rect 52395 18283 52437 18292
rect 52587 18332 52629 18341
rect 52587 18292 52588 18332
rect 52628 18292 52629 18332
rect 52587 18283 52629 18292
rect 576 18164 52800 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 52800 18164
rect 576 18100 52800 18124
rect 8619 17996 8661 18005
rect 8619 17956 8620 17996
rect 8660 17956 8661 17996
rect 8619 17947 8661 17956
rect 22443 17996 22485 18005
rect 22443 17956 22444 17996
rect 22484 17956 22485 17996
rect 22443 17947 22485 17956
rect 26475 17996 26517 18005
rect 26475 17956 26476 17996
rect 26516 17956 26517 17996
rect 26475 17947 26517 17956
rect 33387 17996 33429 18005
rect 33387 17956 33388 17996
rect 33428 17956 33429 17996
rect 33387 17947 33429 17956
rect 36459 17996 36501 18005
rect 36459 17956 36460 17996
rect 36500 17956 36501 17996
rect 36459 17947 36501 17956
rect 46347 17996 46389 18005
rect 46347 17956 46348 17996
rect 46388 17956 46389 17996
rect 46347 17947 46389 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 8323 17912 8381 17913
rect 8323 17872 8332 17912
rect 8372 17872 8381 17912
rect 8323 17871 8381 17872
rect 26755 17912 26813 17913
rect 26755 17872 26764 17912
rect 26804 17872 26813 17912
rect 26755 17871 26813 17872
rect 27723 17912 27765 17921
rect 27723 17872 27724 17912
rect 27764 17872 27765 17912
rect 27723 17863 27765 17872
rect 34731 17912 34773 17921
rect 34731 17872 34732 17912
rect 34772 17872 34773 17912
rect 34731 17863 34773 17872
rect 36747 17912 36789 17921
rect 36747 17872 36748 17912
rect 36788 17872 36789 17912
rect 36747 17863 36789 17872
rect 37803 17912 37845 17921
rect 37803 17872 37804 17912
rect 37844 17872 37845 17912
rect 37803 17863 37845 17872
rect 48459 17912 48501 17921
rect 48459 17872 48460 17912
rect 48500 17872 48501 17912
rect 48459 17863 48501 17872
rect 50091 17912 50133 17921
rect 50091 17872 50092 17912
rect 50132 17872 50133 17912
rect 50091 17863 50133 17872
rect 1699 17828 1757 17829
rect 1699 17788 1708 17828
rect 1748 17788 1757 17828
rect 1699 17787 1757 17788
rect 22243 17828 22301 17829
rect 22243 17788 22252 17828
rect 22292 17788 22301 17828
rect 22243 17787 22301 17788
rect 46531 17828 46589 17829
rect 46531 17788 46540 17828
rect 46580 17788 46589 17828
rect 46531 17787 46589 17788
rect 48259 17828 48317 17829
rect 48259 17788 48268 17828
rect 48308 17788 48317 17828
rect 48259 17787 48317 17788
rect 49411 17828 49469 17829
rect 49411 17788 49420 17828
rect 49460 17788 49469 17828
rect 49411 17787 49469 17788
rect 49891 17758 49949 17759
rect 7651 17744 7709 17745
rect 7651 17704 7660 17744
rect 7700 17704 7709 17744
rect 7651 17703 7709 17704
rect 7947 17744 7989 17753
rect 7947 17704 7948 17744
rect 7988 17704 7989 17744
rect 7947 17695 7989 17704
rect 8523 17744 8565 17753
rect 8523 17704 8524 17744
rect 8564 17704 8565 17744
rect 8523 17695 8565 17704
rect 8707 17744 8765 17745
rect 8707 17704 8716 17744
rect 8756 17704 8765 17744
rect 8707 17703 8765 17704
rect 22635 17744 22677 17753
rect 22635 17704 22636 17744
rect 22676 17704 22677 17744
rect 22635 17695 22677 17704
rect 22827 17744 22869 17753
rect 22827 17704 22828 17744
rect 22868 17704 22869 17744
rect 22827 17695 22869 17704
rect 22915 17744 22973 17745
rect 22915 17704 22924 17744
rect 22964 17704 22973 17744
rect 22915 17703 22973 17704
rect 23491 17744 23549 17745
rect 23491 17704 23500 17744
rect 23540 17704 23549 17744
rect 23491 17703 23549 17704
rect 24355 17744 24413 17745
rect 24355 17704 24364 17744
rect 24404 17704 24413 17744
rect 24355 17703 24413 17704
rect 26371 17744 26429 17745
rect 26371 17704 26380 17744
rect 26420 17704 26429 17744
rect 26371 17703 26429 17704
rect 26571 17744 26613 17753
rect 26571 17704 26572 17744
rect 26612 17704 26613 17744
rect 26571 17695 26613 17704
rect 27051 17744 27093 17753
rect 27051 17704 27052 17744
rect 27092 17704 27093 17744
rect 27051 17695 27093 17704
rect 27147 17744 27189 17753
rect 27147 17704 27148 17744
rect 27188 17704 27189 17744
rect 27147 17695 27189 17704
rect 27427 17744 27485 17745
rect 27427 17704 27436 17744
rect 27476 17704 27485 17744
rect 27427 17703 27485 17704
rect 29931 17744 29973 17753
rect 29931 17704 29932 17744
rect 29972 17704 29973 17744
rect 29931 17695 29973 17704
rect 30123 17744 30165 17753
rect 30123 17704 30124 17744
rect 30164 17704 30165 17744
rect 30123 17695 30165 17704
rect 30211 17744 30269 17745
rect 30211 17704 30220 17744
rect 30260 17704 30269 17744
rect 30211 17703 30269 17704
rect 30787 17744 30845 17745
rect 30787 17704 30796 17744
rect 30836 17704 30845 17744
rect 30787 17703 30845 17704
rect 31651 17744 31709 17745
rect 31651 17704 31660 17744
rect 31700 17704 31709 17744
rect 31651 17703 31709 17704
rect 33283 17744 33341 17745
rect 33283 17704 33292 17744
rect 33332 17704 33341 17744
rect 33283 17703 33341 17704
rect 33483 17744 33525 17753
rect 33483 17704 33484 17744
rect 33524 17704 33525 17744
rect 33483 17695 33525 17704
rect 34147 17744 34205 17745
rect 34147 17704 34156 17744
rect 34196 17704 34205 17744
rect 34147 17703 34205 17704
rect 34347 17744 34389 17753
rect 34347 17704 34348 17744
rect 34388 17704 34389 17744
rect 34347 17695 34389 17704
rect 36355 17744 36413 17745
rect 36355 17704 36364 17744
rect 36404 17704 36413 17744
rect 36355 17703 36413 17704
rect 36555 17744 36597 17753
rect 36555 17704 36556 17744
rect 36596 17704 36597 17744
rect 36555 17695 36597 17704
rect 39819 17744 39861 17753
rect 39819 17704 39820 17744
rect 39860 17704 39861 17744
rect 39819 17695 39861 17704
rect 40195 17744 40253 17745
rect 40195 17704 40204 17744
rect 40244 17704 40253 17744
rect 40195 17703 40253 17704
rect 41059 17744 41117 17745
rect 41059 17704 41068 17744
rect 41108 17704 41117 17744
rect 41059 17703 41117 17704
rect 42699 17744 42741 17753
rect 42699 17704 42700 17744
rect 42740 17704 42741 17744
rect 42699 17695 42741 17704
rect 42891 17744 42933 17753
rect 42891 17704 42892 17744
rect 42932 17704 42933 17744
rect 42891 17695 42933 17704
rect 42979 17744 43037 17745
rect 42979 17704 42988 17744
rect 43028 17704 43037 17744
rect 42979 17703 43037 17704
rect 43555 17744 43613 17745
rect 43555 17704 43564 17744
rect 43604 17704 43613 17744
rect 43555 17703 43613 17704
rect 44419 17744 44477 17745
rect 44419 17704 44428 17744
rect 44468 17704 44477 17744
rect 44419 17703 44477 17704
rect 46051 17744 46109 17745
rect 46051 17704 46060 17744
rect 46100 17704 46109 17744
rect 46051 17703 46109 17704
rect 46155 17744 46197 17753
rect 46155 17704 46156 17744
rect 46196 17704 46197 17744
rect 46155 17695 46197 17704
rect 46347 17744 46389 17753
rect 46347 17704 46348 17744
rect 46388 17704 46389 17744
rect 46347 17695 46389 17704
rect 48643 17744 48701 17745
rect 48643 17704 48652 17744
rect 48692 17704 48701 17744
rect 48643 17703 48701 17704
rect 48747 17744 48789 17753
rect 48747 17704 48748 17744
rect 48788 17704 48789 17744
rect 48747 17695 48789 17704
rect 48939 17744 48981 17753
rect 48939 17704 48940 17744
rect 48980 17704 48981 17744
rect 48939 17695 48981 17704
rect 49795 17744 49853 17745
rect 49795 17704 49804 17744
rect 49844 17704 49853 17744
rect 49891 17718 49900 17758
rect 49940 17718 49949 17758
rect 49891 17717 49949 17718
rect 50091 17744 50133 17753
rect 49795 17703 49853 17704
rect 50091 17704 50092 17744
rect 50132 17704 50133 17744
rect 50091 17695 50133 17704
rect 50283 17744 50325 17753
rect 50283 17704 50284 17744
rect 50324 17704 50325 17744
rect 50283 17695 50325 17704
rect 50659 17744 50717 17745
rect 50659 17704 50668 17744
rect 50708 17704 50717 17744
rect 50659 17703 50717 17704
rect 51523 17744 51581 17745
rect 51523 17704 51532 17744
rect 51572 17704 51581 17744
rect 51523 17703 51581 17704
rect 8043 17660 8085 17669
rect 8043 17620 8044 17660
rect 8084 17620 8085 17660
rect 8043 17611 8085 17620
rect 22731 17660 22773 17669
rect 22731 17620 22732 17660
rect 22772 17620 22773 17660
rect 22731 17611 22773 17620
rect 23115 17660 23157 17669
rect 23115 17620 23116 17660
rect 23156 17620 23157 17660
rect 23115 17611 23157 17620
rect 30027 17660 30069 17669
rect 30027 17620 30028 17660
rect 30068 17620 30069 17660
rect 30027 17611 30069 17620
rect 30411 17660 30453 17669
rect 30411 17620 30412 17660
rect 30452 17620 30453 17660
rect 30411 17611 30453 17620
rect 34251 17660 34293 17669
rect 34251 17620 34252 17660
rect 34292 17620 34293 17660
rect 34251 17611 34293 17620
rect 42795 17660 42837 17669
rect 42795 17620 42796 17660
rect 42836 17620 42837 17660
rect 42795 17611 42837 17620
rect 43179 17660 43221 17669
rect 43179 17620 43180 17660
rect 43220 17620 43221 17660
rect 43179 17611 43221 17620
rect 1515 17576 1557 17585
rect 1515 17536 1516 17576
rect 1556 17536 1557 17576
rect 1515 17527 1557 17536
rect 25507 17576 25565 17577
rect 25507 17536 25516 17576
rect 25556 17536 25565 17576
rect 25507 17535 25565 17536
rect 32803 17576 32861 17577
rect 32803 17536 32812 17576
rect 32852 17536 32861 17576
rect 32803 17535 32861 17536
rect 42211 17576 42269 17577
rect 42211 17536 42220 17576
rect 42260 17536 42269 17576
rect 42211 17535 42269 17536
rect 45571 17576 45629 17577
rect 45571 17536 45580 17576
rect 45620 17536 45629 17576
rect 45571 17535 45629 17536
rect 46731 17576 46773 17585
rect 46731 17536 46732 17576
rect 46772 17536 46773 17576
rect 46731 17527 46773 17536
rect 48835 17576 48893 17577
rect 48835 17536 48844 17576
rect 48884 17536 48893 17576
rect 48835 17535 48893 17536
rect 49611 17576 49653 17585
rect 49611 17536 49612 17576
rect 49652 17536 49653 17576
rect 49611 17527 49653 17536
rect 52675 17576 52733 17577
rect 52675 17536 52684 17576
rect 52724 17536 52733 17576
rect 52675 17535 52733 17536
rect 576 17408 52800 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 52800 17408
rect 576 17344 52800 17368
rect 2475 17240 2517 17249
rect 2475 17200 2476 17240
rect 2516 17200 2517 17240
rect 2475 17191 2517 17200
rect 26851 17240 26909 17241
rect 26851 17200 26860 17240
rect 26900 17200 26909 17240
rect 26851 17199 26909 17200
rect 41635 17240 41693 17241
rect 41635 17200 41644 17240
rect 41684 17200 41693 17240
rect 41635 17199 41693 17200
rect 22827 17156 22869 17165
rect 22827 17116 22828 17156
rect 22868 17116 22869 17156
rect 22827 17107 22869 17116
rect 23211 17156 23253 17165
rect 23211 17116 23212 17156
rect 23252 17116 23253 17156
rect 23211 17107 23253 17116
rect 27243 17156 27285 17165
rect 27243 17116 27244 17156
rect 27284 17116 27285 17156
rect 27243 17107 27285 17116
rect 33867 17156 33909 17165
rect 33867 17116 33868 17156
rect 33908 17116 33909 17156
rect 33867 17107 33909 17116
rect 44139 17156 44181 17165
rect 44139 17116 44140 17156
rect 44180 17116 44181 17156
rect 44139 17107 44181 17116
rect 45771 17156 45813 17165
rect 45771 17116 45772 17156
rect 45812 17116 45813 17156
rect 45771 17107 45813 17116
rect 51339 17156 51381 17165
rect 51339 17116 51340 17156
rect 51380 17116 51381 17156
rect 51339 17107 51381 17116
rect 22731 17072 22773 17081
rect 22731 17032 22732 17072
rect 22772 17032 22773 17072
rect 22731 17023 22773 17032
rect 22915 17072 22973 17073
rect 22915 17032 22924 17072
rect 22964 17032 22973 17072
rect 22915 17031 22973 17032
rect 23107 17072 23165 17073
rect 23107 17032 23116 17072
rect 23156 17032 23165 17072
rect 23107 17031 23165 17032
rect 23307 17072 23349 17081
rect 23307 17032 23308 17072
rect 23348 17032 23349 17072
rect 23307 17023 23349 17032
rect 26763 17072 26805 17081
rect 26763 17032 26764 17072
rect 26804 17032 26805 17072
rect 26763 17023 26805 17032
rect 26955 17072 26997 17081
rect 26955 17032 26956 17072
rect 26996 17032 26997 17072
rect 26955 17023 26997 17032
rect 27043 17072 27101 17073
rect 27043 17032 27052 17072
rect 27092 17032 27101 17072
rect 27043 17031 27101 17032
rect 27619 17072 27677 17073
rect 27619 17032 27628 17072
rect 27668 17032 27677 17072
rect 27619 17031 27677 17032
rect 28483 17072 28541 17073
rect 28483 17032 28492 17072
rect 28532 17032 28541 17072
rect 28483 17031 28541 17032
rect 30507 17072 30549 17081
rect 30507 17032 30508 17072
rect 30548 17032 30549 17072
rect 30507 17023 30549 17032
rect 30691 17072 30749 17073
rect 30691 17032 30700 17072
rect 30740 17032 30749 17072
rect 30691 17031 30749 17032
rect 33771 17072 33813 17081
rect 33771 17032 33772 17072
rect 33812 17032 33813 17072
rect 33771 17023 33813 17032
rect 33963 17072 34005 17081
rect 33963 17032 33964 17072
rect 34004 17032 34005 17072
rect 33963 17023 34005 17032
rect 34051 17072 34109 17073
rect 34051 17032 34060 17072
rect 34100 17032 34109 17072
rect 34051 17031 34109 17032
rect 34251 17072 34293 17081
rect 34251 17032 34252 17072
rect 34292 17032 34293 17072
rect 34251 17023 34293 17032
rect 34627 17072 34685 17073
rect 34627 17032 34636 17072
rect 34676 17032 34685 17072
rect 34627 17031 34685 17032
rect 35491 17072 35549 17073
rect 35491 17032 35500 17072
rect 35540 17032 35549 17072
rect 35491 17031 35549 17032
rect 36931 17072 36989 17073
rect 36931 17032 36940 17072
rect 36980 17032 36989 17072
rect 36931 17031 36989 17032
rect 37131 17072 37173 17081
rect 37131 17032 37132 17072
rect 37172 17032 37173 17072
rect 37131 17023 37173 17032
rect 37323 17072 37365 17081
rect 37323 17032 37324 17072
rect 37364 17032 37365 17072
rect 37323 17023 37365 17032
rect 37699 17072 37757 17073
rect 37699 17032 37708 17072
rect 37748 17032 37757 17072
rect 37699 17031 37757 17032
rect 38563 17072 38621 17073
rect 38563 17032 38572 17072
rect 38612 17032 38621 17072
rect 38563 17031 38621 17032
rect 41739 17072 41781 17081
rect 41739 17032 41740 17072
rect 41780 17032 41781 17072
rect 41739 17023 41781 17032
rect 41835 17072 41877 17081
rect 41835 17032 41836 17072
rect 41876 17032 41877 17072
rect 41835 17023 41877 17032
rect 41931 17072 41973 17081
rect 41931 17032 41932 17072
rect 41972 17032 41973 17072
rect 41931 17023 41973 17032
rect 42211 17072 42269 17073
rect 42211 17032 42220 17072
rect 42260 17032 42269 17072
rect 42211 17031 42269 17032
rect 42507 17072 42549 17081
rect 42507 17032 42508 17072
rect 42548 17032 42549 17072
rect 42507 17023 42549 17032
rect 42603 17072 42645 17081
rect 42603 17032 42604 17072
rect 42644 17032 42645 17072
rect 42603 17023 42645 17032
rect 44043 17072 44085 17081
rect 44043 17032 44044 17072
rect 44084 17032 44085 17072
rect 44043 17023 44085 17032
rect 44227 17072 44285 17073
rect 44227 17032 44236 17072
rect 44276 17032 44285 17072
rect 44227 17031 44285 17032
rect 45379 17072 45437 17073
rect 45379 17032 45388 17072
rect 45428 17032 45437 17072
rect 45379 17031 45437 17032
rect 45675 17072 45717 17081
rect 45675 17032 45676 17072
rect 45716 17032 45717 17072
rect 45675 17023 45717 17032
rect 46251 17072 46293 17081
rect 46251 17032 46252 17072
rect 46292 17032 46293 17072
rect 46251 17023 46293 17032
rect 46627 17072 46685 17073
rect 46627 17032 46636 17072
rect 46676 17032 46685 17072
rect 46627 17031 46685 17032
rect 47491 17072 47549 17073
rect 47491 17032 47500 17072
rect 47540 17032 47549 17072
rect 47491 17031 47549 17032
rect 49123 17072 49181 17073
rect 49123 17032 49132 17072
rect 49172 17032 49181 17072
rect 49123 17031 49181 17032
rect 49227 17072 49269 17081
rect 49227 17032 49228 17072
rect 49268 17032 49269 17072
rect 49227 17023 49269 17032
rect 49419 17072 49461 17081
rect 49419 17032 49420 17072
rect 49460 17032 49461 17072
rect 49419 17023 49461 17032
rect 50371 17072 50429 17073
rect 50371 17032 50380 17072
rect 50420 17032 50429 17072
rect 50371 17031 50429 17032
rect 50667 17072 50709 17081
rect 50667 17032 50668 17072
rect 50708 17032 50709 17072
rect 50667 17023 50709 17032
rect 50763 17072 50805 17081
rect 50763 17032 50764 17072
rect 50804 17032 50805 17072
rect 50763 17023 50805 17032
rect 51235 17072 51293 17073
rect 51235 17032 51244 17072
rect 51284 17032 51293 17072
rect 51235 17031 51293 17032
rect 51435 17072 51477 17081
rect 51435 17032 51436 17072
rect 51476 17032 51477 17072
rect 51435 17023 51477 17032
rect 52291 17072 52349 17073
rect 52291 17032 52300 17072
rect 52340 17032 52349 17072
rect 52291 17031 52349 17032
rect 52579 17072 52637 17073
rect 52579 17032 52588 17072
rect 52628 17032 52637 17072
rect 52579 17031 52637 17032
rect 51619 17001 51677 17002
rect 2659 16988 2717 16989
rect 2659 16948 2668 16988
rect 2708 16948 2717 16988
rect 2659 16947 2717 16948
rect 33379 16988 33437 16989
rect 33379 16948 33388 16988
rect 33428 16948 33437 16988
rect 33379 16947 33437 16948
rect 41059 16988 41117 16989
rect 41059 16948 41068 16988
rect 41108 16948 41117 16988
rect 41059 16947 41117 16948
rect 41443 16988 41501 16989
rect 41443 16948 41452 16988
rect 41492 16948 41501 16988
rect 41443 16947 41501 16948
rect 43075 16988 43133 16989
rect 43075 16948 43084 16988
rect 43124 16948 43133 16988
rect 43075 16947 43133 16948
rect 44515 16988 44573 16989
rect 44515 16948 44524 16988
rect 44564 16948 44573 16988
rect 44515 16947 44573 16948
rect 44899 16988 44957 16989
rect 44899 16948 44908 16988
rect 44948 16948 44957 16988
rect 44899 16947 44957 16948
rect 48651 16988 48693 16997
rect 48651 16948 48652 16988
rect 48692 16948 48693 16988
rect 48651 16939 48693 16948
rect 49891 16988 49949 16989
rect 49891 16948 49900 16988
rect 49940 16948 49949 16988
rect 51619 16961 51628 17001
rect 51668 16961 51677 17001
rect 51619 16960 51677 16961
rect 52395 16988 52437 16997
rect 49891 16947 49949 16948
rect 52395 16948 52396 16988
rect 52436 16948 52437 16988
rect 52395 16939 52437 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 23691 16904 23733 16913
rect 23691 16864 23692 16904
rect 23732 16864 23733 16904
rect 23691 16855 23733 16864
rect 30603 16904 30645 16913
rect 30603 16864 30604 16904
rect 30644 16864 30645 16904
rect 30603 16855 30645 16864
rect 30891 16904 30933 16913
rect 30891 16864 30892 16904
rect 30932 16864 30933 16904
rect 30891 16855 30933 16864
rect 36643 16904 36701 16905
rect 36643 16864 36652 16904
rect 36692 16864 36701 16904
rect 36643 16863 36701 16864
rect 40875 16904 40917 16913
rect 40875 16864 40876 16904
rect 40916 16864 40917 16904
rect 40875 16855 40917 16864
rect 42883 16904 42941 16905
rect 42883 16864 42892 16904
rect 42932 16864 42941 16904
rect 42883 16863 42941 16864
rect 43659 16904 43701 16913
rect 43659 16864 43660 16904
rect 43700 16864 43701 16904
rect 43659 16855 43701 16864
rect 44715 16904 44757 16913
rect 44715 16864 44716 16904
rect 44756 16864 44757 16904
rect 44715 16855 44757 16864
rect 52683 16904 52725 16913
rect 52683 16864 52684 16904
rect 52724 16864 52725 16904
rect 52683 16855 52725 16864
rect 29635 16820 29693 16821
rect 29635 16780 29644 16820
rect 29684 16780 29693 16820
rect 29635 16779 29693 16780
rect 33579 16820 33621 16829
rect 33579 16780 33580 16820
rect 33620 16780 33621 16820
rect 33579 16771 33621 16780
rect 37035 16820 37077 16829
rect 37035 16780 37036 16820
rect 37076 16780 37077 16820
rect 37035 16771 37077 16780
rect 39715 16820 39773 16821
rect 39715 16780 39724 16820
rect 39764 16780 39773 16820
rect 39715 16779 39773 16780
rect 41259 16820 41301 16829
rect 41259 16780 41260 16820
rect 41300 16780 41301 16820
rect 41259 16771 41301 16780
rect 43275 16820 43317 16829
rect 43275 16780 43276 16820
rect 43316 16780 43317 16820
rect 43275 16771 43317 16780
rect 45099 16820 45141 16829
rect 45099 16780 45100 16820
rect 45140 16780 45141 16820
rect 45099 16771 45141 16780
rect 46051 16820 46109 16821
rect 46051 16780 46060 16820
rect 46100 16780 46109 16820
rect 46051 16779 46109 16780
rect 49419 16820 49461 16829
rect 49419 16780 49420 16820
rect 49460 16780 49461 16820
rect 49419 16771 49461 16780
rect 50091 16820 50133 16829
rect 50091 16780 50092 16820
rect 50132 16780 50133 16820
rect 50091 16771 50133 16780
rect 51043 16820 51101 16821
rect 51043 16780 51052 16820
rect 51092 16780 51101 16820
rect 51043 16779 51101 16780
rect 51819 16820 51861 16829
rect 51819 16780 51820 16820
rect 51860 16780 51861 16820
rect 51819 16771 51861 16780
rect 576 16652 79584 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 79584 16652
rect 576 16588 79584 16612
rect 4203 16484 4245 16493
rect 4203 16444 4204 16484
rect 4244 16444 4245 16484
rect 4203 16435 4245 16444
rect 34635 16484 34677 16493
rect 34635 16444 34636 16484
rect 34676 16444 34677 16484
rect 34635 16435 34677 16444
rect 37995 16484 38037 16493
rect 37995 16444 37996 16484
rect 38036 16444 38037 16484
rect 37995 16435 38037 16444
rect 42691 16484 42749 16485
rect 42691 16444 42700 16484
rect 42740 16444 42749 16484
rect 42691 16443 42749 16444
rect 42987 16484 43029 16493
rect 42987 16444 42988 16484
rect 43028 16444 43029 16484
rect 42987 16435 43029 16444
rect 45667 16484 45725 16485
rect 45667 16444 45676 16484
rect 45716 16444 45725 16484
rect 45667 16443 45725 16444
rect 45963 16484 46005 16493
rect 45963 16444 45964 16484
rect 46004 16444 46005 16484
rect 45963 16435 46005 16444
rect 51339 16484 51381 16493
rect 51339 16444 51340 16484
rect 51380 16444 51381 16484
rect 51339 16435 51381 16444
rect 54507 16484 54549 16493
rect 54507 16444 54508 16484
rect 54548 16444 54549 16484
rect 54507 16435 54549 16444
rect 54891 16484 54933 16493
rect 54891 16444 54892 16484
rect 54932 16444 54933 16484
rect 54891 16435 54933 16444
rect 55755 16484 55797 16493
rect 55755 16444 55756 16484
rect 55796 16444 55797 16484
rect 55755 16435 55797 16444
rect 56235 16484 56277 16493
rect 56235 16444 56236 16484
rect 56276 16444 56277 16484
rect 56235 16435 56277 16444
rect 56619 16484 56661 16493
rect 56619 16444 56620 16484
rect 56660 16444 56661 16484
rect 56619 16435 56661 16444
rect 57387 16484 57429 16493
rect 57387 16444 57388 16484
rect 57428 16444 57429 16484
rect 57387 16435 57429 16444
rect 58059 16484 58101 16493
rect 58059 16444 58060 16484
rect 58100 16444 58101 16484
rect 58059 16435 58101 16444
rect 58347 16484 58389 16493
rect 58347 16444 58348 16484
rect 58388 16444 58389 16484
rect 58347 16435 58389 16444
rect 58635 16484 58677 16493
rect 58635 16444 58636 16484
rect 58676 16444 58677 16484
rect 58635 16435 58677 16444
rect 60171 16484 60213 16493
rect 60171 16444 60172 16484
rect 60212 16444 60213 16484
rect 60171 16435 60213 16444
rect 60651 16484 60693 16493
rect 60651 16444 60652 16484
rect 60692 16444 60693 16484
rect 60651 16435 60693 16444
rect 61515 16484 61557 16493
rect 61515 16444 61516 16484
rect 61556 16444 61557 16484
rect 61515 16435 61557 16444
rect 62187 16484 62229 16493
rect 62187 16444 62188 16484
rect 62228 16444 62229 16484
rect 62187 16435 62229 16444
rect 62475 16484 62517 16493
rect 62475 16444 62476 16484
rect 62516 16444 62517 16484
rect 62475 16435 62517 16444
rect 63051 16484 63093 16493
rect 63051 16444 63052 16484
rect 63092 16444 63093 16484
rect 63051 16435 63093 16444
rect 63339 16484 63381 16493
rect 63339 16444 63340 16484
rect 63380 16444 63381 16484
rect 63339 16435 63381 16444
rect 63627 16484 63669 16493
rect 63627 16444 63628 16484
rect 63668 16444 63669 16484
rect 63627 16435 63669 16444
rect 63915 16484 63957 16493
rect 63915 16444 63916 16484
rect 63956 16444 63957 16484
rect 63915 16435 63957 16444
rect 64587 16484 64629 16493
rect 64587 16444 64588 16484
rect 64628 16444 64629 16484
rect 64587 16435 64629 16444
rect 65067 16484 65109 16493
rect 65067 16444 65068 16484
rect 65108 16444 65109 16484
rect 65067 16435 65109 16444
rect 65451 16484 65493 16493
rect 65451 16444 65452 16484
rect 65492 16444 65493 16484
rect 65451 16435 65493 16444
rect 65835 16484 65877 16493
rect 65835 16444 65836 16484
rect 65876 16444 65877 16484
rect 65835 16435 65877 16444
rect 66603 16484 66645 16493
rect 66603 16444 66604 16484
rect 66644 16444 66645 16484
rect 66603 16435 66645 16444
rect 67083 16484 67125 16493
rect 67083 16444 67084 16484
rect 67124 16444 67125 16484
rect 67083 16435 67125 16444
rect 67467 16484 67509 16493
rect 67467 16444 67468 16484
rect 67508 16444 67509 16484
rect 67467 16435 67509 16444
rect 67851 16484 67893 16493
rect 67851 16444 67852 16484
rect 67892 16444 67893 16484
rect 67851 16435 67893 16444
rect 68235 16484 68277 16493
rect 68235 16444 68236 16484
rect 68276 16444 68277 16484
rect 68235 16435 68277 16444
rect 69099 16484 69141 16493
rect 69099 16444 69100 16484
rect 69140 16444 69141 16484
rect 69099 16435 69141 16444
rect 69483 16484 69525 16493
rect 69483 16444 69484 16484
rect 69524 16444 69525 16484
rect 69483 16435 69525 16444
rect 69867 16484 69909 16493
rect 69867 16444 69868 16484
rect 69908 16444 69909 16484
rect 69867 16435 69909 16444
rect 70251 16484 70293 16493
rect 70251 16444 70252 16484
rect 70292 16444 70293 16484
rect 70251 16435 70293 16444
rect 70635 16484 70677 16493
rect 70635 16444 70636 16484
rect 70676 16444 70677 16484
rect 70635 16435 70677 16444
rect 71019 16484 71061 16493
rect 71019 16444 71020 16484
rect 71060 16444 71061 16484
rect 71019 16435 71061 16444
rect 71403 16484 71445 16493
rect 71403 16444 71404 16484
rect 71444 16444 71445 16484
rect 71403 16435 71445 16444
rect 71883 16484 71925 16493
rect 71883 16444 71884 16484
rect 71924 16444 71925 16484
rect 71883 16435 71925 16444
rect 72267 16484 72309 16493
rect 72267 16444 72268 16484
rect 72308 16444 72309 16484
rect 72267 16435 72309 16444
rect 72651 16484 72693 16493
rect 72651 16444 72652 16484
rect 72692 16444 72693 16484
rect 72651 16435 72693 16444
rect 73035 16484 73077 16493
rect 73035 16444 73036 16484
rect 73076 16444 73077 16484
rect 73035 16435 73077 16444
rect 73419 16484 73461 16493
rect 73419 16444 73420 16484
rect 73460 16444 73461 16484
rect 73419 16435 73461 16444
rect 74283 16484 74325 16493
rect 74283 16444 74284 16484
rect 74324 16444 74325 16484
rect 74283 16435 74325 16444
rect 74667 16484 74709 16493
rect 74667 16444 74668 16484
rect 74708 16444 74709 16484
rect 74667 16435 74709 16444
rect 75051 16484 75093 16493
rect 75051 16444 75052 16484
rect 75092 16444 75093 16484
rect 75051 16435 75093 16444
rect 75435 16484 75477 16493
rect 75435 16444 75436 16484
rect 75476 16444 75477 16484
rect 75435 16435 75477 16444
rect 75819 16484 75861 16493
rect 75819 16444 75820 16484
rect 75860 16444 75861 16484
rect 75819 16435 75861 16444
rect 76491 16484 76533 16493
rect 76491 16444 76492 16484
rect 76532 16444 76533 16484
rect 76491 16435 76533 16444
rect 76875 16484 76917 16493
rect 76875 16444 76876 16484
rect 76916 16444 76917 16484
rect 76875 16435 76917 16444
rect 77259 16484 77301 16493
rect 77259 16444 77260 16484
rect 77300 16444 77301 16484
rect 77259 16435 77301 16444
rect 77547 16484 77589 16493
rect 77547 16444 77548 16484
rect 77588 16444 77589 16484
rect 77547 16435 77589 16444
rect 77931 16484 77973 16493
rect 77931 16444 77932 16484
rect 77972 16444 77973 16484
rect 77931 16435 77973 16444
rect 78315 16484 78357 16493
rect 78315 16444 78316 16484
rect 78356 16444 78357 16484
rect 78315 16435 78357 16444
rect 78699 16484 78741 16493
rect 78699 16444 78700 16484
rect 78740 16444 78741 16484
rect 78699 16435 78741 16444
rect 78987 16484 79029 16493
rect 78987 16444 78988 16484
rect 79028 16444 79029 16484
rect 78987 16435 79029 16444
rect 79275 16484 79317 16493
rect 79275 16444 79276 16484
rect 79316 16444 79317 16484
rect 79275 16435 79317 16444
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 1515 16400 1557 16409
rect 1515 16360 1516 16400
rect 1556 16360 1557 16400
rect 1515 16351 1557 16360
rect 2379 16400 2421 16409
rect 2379 16360 2380 16400
rect 2420 16360 2421 16400
rect 2379 16351 2421 16360
rect 34339 16400 34397 16401
rect 34339 16360 34348 16400
rect 34388 16360 34397 16400
rect 34339 16359 34397 16360
rect 36739 16400 36797 16401
rect 36739 16360 36748 16400
rect 36788 16360 36797 16400
rect 36739 16359 36797 16360
rect 46827 16400 46869 16409
rect 46827 16360 46828 16400
rect 46868 16360 46869 16400
rect 46827 16351 46869 16360
rect 53163 16400 53205 16409
rect 53163 16360 53164 16400
rect 53204 16360 53205 16400
rect 53163 16351 53205 16360
rect 53643 16400 53685 16409
rect 53643 16360 53644 16400
rect 53684 16360 53685 16400
rect 53643 16351 53685 16360
rect 57579 16400 57621 16409
rect 57579 16360 57580 16400
rect 57620 16360 57621 16400
rect 57579 16351 57621 16360
rect 61035 16400 61077 16409
rect 61035 16360 61036 16400
rect 61076 16360 61077 16400
rect 61035 16351 61077 16360
rect 1987 16316 2045 16317
rect 1987 16276 1996 16316
rect 2036 16276 2045 16316
rect 1987 16275 2045 16276
rect 2563 16316 2621 16317
rect 2563 16276 2572 16316
rect 2612 16276 2621 16316
rect 2563 16275 2621 16276
rect 2755 16316 2813 16317
rect 2755 16276 2764 16316
rect 2804 16276 2813 16316
rect 2755 16275 2813 16276
rect 4387 16316 4445 16317
rect 4387 16276 4396 16316
rect 4436 16276 4445 16316
rect 4387 16275 4445 16276
rect 46627 16316 46685 16317
rect 46627 16276 46636 16316
rect 46676 16276 46685 16316
rect 46627 16275 46685 16276
rect 61699 16316 61757 16317
rect 61699 16276 61708 16316
rect 61748 16276 61757 16316
rect 61699 16275 61757 16276
rect 27352 16247 27394 16256
rect 3339 16232 3381 16241
rect 3339 16192 3340 16232
rect 3380 16192 3381 16232
rect 3339 16183 3381 16192
rect 3523 16232 3581 16233
rect 3523 16192 3532 16232
rect 3572 16192 3581 16232
rect 3523 16191 3581 16192
rect 4963 16232 5021 16233
rect 4963 16192 4972 16232
rect 5012 16192 5021 16232
rect 4963 16191 5021 16192
rect 5827 16232 5885 16233
rect 5827 16192 5836 16232
rect 5876 16192 5885 16232
rect 27352 16207 27353 16247
rect 27393 16207 27394 16247
rect 27352 16198 27394 16207
rect 27531 16232 27573 16241
rect 5827 16191 5885 16192
rect 27531 16192 27532 16232
rect 27572 16192 27573 16232
rect 27531 16183 27573 16192
rect 31363 16232 31421 16233
rect 31363 16192 31372 16232
rect 31412 16192 31421 16232
rect 31363 16191 31421 16192
rect 32227 16232 32285 16233
rect 32227 16192 32236 16232
rect 32276 16192 32285 16232
rect 32227 16191 32285 16192
rect 33667 16232 33725 16233
rect 33667 16192 33676 16232
rect 33716 16192 33725 16232
rect 33667 16191 33725 16192
rect 33963 16232 34005 16241
rect 33963 16192 33964 16232
rect 34004 16192 34005 16232
rect 33963 16183 34005 16192
rect 34539 16232 34581 16241
rect 34539 16192 34540 16232
rect 34580 16192 34581 16232
rect 34539 16183 34581 16192
rect 34723 16232 34781 16233
rect 34723 16192 34732 16232
rect 34772 16192 34781 16232
rect 34723 16191 34781 16192
rect 36355 16232 36413 16233
rect 36355 16192 36364 16232
rect 36404 16192 36413 16232
rect 36355 16191 36413 16192
rect 36459 16232 36501 16241
rect 36459 16192 36460 16232
rect 36500 16192 36501 16232
rect 36459 16183 36501 16192
rect 36555 16232 36597 16241
rect 36555 16192 36556 16232
rect 36596 16192 36597 16232
rect 36555 16183 36597 16192
rect 37131 16232 37173 16241
rect 37131 16192 37132 16232
rect 37172 16192 37173 16232
rect 37131 16183 37173 16192
rect 37411 16232 37469 16233
rect 37411 16192 37420 16232
rect 37460 16192 37469 16232
rect 37411 16191 37469 16192
rect 37699 16232 37757 16233
rect 37699 16192 37708 16232
rect 37748 16192 37757 16232
rect 37699 16191 37757 16192
rect 37803 16232 37845 16241
rect 37803 16192 37804 16232
rect 37844 16192 37845 16232
rect 37803 16183 37845 16192
rect 37995 16232 38037 16241
rect 37995 16192 37996 16232
rect 38036 16192 38037 16232
rect 37995 16183 38037 16192
rect 39915 16232 39957 16241
rect 39915 16192 39916 16232
rect 39956 16192 39957 16232
rect 39915 16183 39957 16192
rect 40099 16232 40157 16233
rect 40099 16192 40108 16232
rect 40148 16192 40157 16232
rect 40099 16191 40157 16192
rect 40675 16232 40733 16233
rect 40675 16192 40684 16232
rect 40724 16192 40733 16232
rect 40675 16191 40733 16192
rect 41539 16232 41597 16233
rect 41539 16192 41548 16232
rect 41588 16192 41597 16232
rect 41539 16191 41597 16192
rect 42891 16232 42933 16241
rect 42891 16192 42892 16232
rect 42932 16192 42933 16232
rect 42891 16183 42933 16192
rect 43075 16232 43133 16233
rect 43075 16192 43084 16232
rect 43124 16192 43133 16232
rect 43075 16191 43133 16192
rect 43651 16232 43709 16233
rect 43651 16192 43660 16232
rect 43700 16192 43709 16232
rect 43651 16191 43709 16192
rect 44515 16232 44573 16233
rect 44515 16192 44524 16232
rect 44564 16192 44573 16232
rect 44515 16191 44573 16192
rect 45963 16232 46005 16241
rect 45963 16192 45964 16232
rect 46004 16192 46005 16232
rect 45963 16183 46005 16192
rect 46155 16232 46197 16241
rect 46155 16192 46156 16232
rect 46196 16192 46197 16232
rect 46155 16183 46197 16192
rect 46243 16232 46301 16233
rect 46243 16192 46252 16232
rect 46292 16192 46301 16232
rect 46243 16191 46301 16192
rect 48651 16232 48693 16241
rect 48651 16192 48652 16232
rect 48692 16192 48693 16232
rect 48651 16183 48693 16192
rect 49027 16232 49085 16233
rect 49027 16192 49036 16232
rect 49076 16192 49085 16232
rect 49027 16191 49085 16192
rect 49891 16232 49949 16233
rect 49891 16192 49900 16232
rect 49940 16192 49949 16232
rect 49891 16191 49949 16192
rect 51243 16232 51285 16241
rect 51243 16192 51244 16232
rect 51284 16192 51285 16232
rect 51243 16183 51285 16192
rect 51427 16232 51485 16233
rect 51427 16192 51436 16232
rect 51476 16192 51485 16232
rect 51427 16191 51485 16192
rect 51619 16232 51677 16233
rect 51619 16192 51628 16232
rect 51668 16192 51677 16232
rect 51619 16191 51677 16192
rect 52587 16232 52629 16241
rect 52587 16192 52588 16232
rect 52628 16192 52629 16232
rect 52587 16183 52629 16192
rect 52779 16232 52821 16241
rect 52779 16192 52780 16232
rect 52820 16192 52821 16232
rect 52779 16183 52821 16192
rect 52867 16232 52925 16233
rect 52867 16192 52876 16232
rect 52916 16192 52925 16232
rect 52867 16191 52925 16192
rect 53059 16232 53117 16233
rect 53059 16192 53068 16232
rect 53108 16192 53117 16232
rect 54403 16232 54461 16233
rect 53059 16191 53117 16192
rect 53268 16219 53310 16228
rect 53268 16179 53269 16219
rect 53309 16179 53310 16219
rect 54403 16192 54412 16232
rect 54452 16192 54461 16232
rect 54403 16191 54461 16192
rect 54787 16232 54845 16233
rect 54787 16192 54796 16232
rect 54836 16192 54845 16232
rect 54787 16191 54845 16192
rect 55267 16232 55325 16233
rect 55267 16192 55276 16232
rect 55316 16192 55325 16232
rect 55267 16191 55325 16192
rect 55651 16232 55709 16233
rect 55651 16192 55660 16232
rect 55700 16192 55709 16232
rect 55651 16191 55709 16192
rect 56131 16232 56189 16233
rect 56131 16192 56140 16232
rect 56180 16192 56189 16232
rect 56131 16191 56189 16192
rect 56515 16232 56573 16233
rect 56515 16192 56524 16232
rect 56564 16192 56573 16232
rect 56515 16191 56573 16192
rect 56899 16232 56957 16233
rect 56899 16192 56908 16232
rect 56948 16192 56957 16232
rect 56899 16191 56957 16192
rect 57283 16232 57341 16233
rect 57283 16192 57292 16232
rect 57332 16192 57341 16232
rect 57283 16191 57341 16192
rect 57955 16232 58013 16233
rect 57955 16192 57964 16232
rect 58004 16192 58013 16232
rect 57955 16191 58013 16192
rect 58243 16232 58301 16233
rect 58243 16192 58252 16232
rect 58292 16192 58301 16232
rect 58243 16191 58301 16192
rect 58531 16232 58589 16233
rect 58531 16192 58540 16232
rect 58580 16192 58589 16232
rect 58531 16191 58589 16192
rect 58915 16232 58973 16233
rect 58915 16192 58924 16232
rect 58964 16192 58973 16232
rect 58915 16191 58973 16192
rect 59299 16232 59357 16233
rect 59299 16192 59308 16232
rect 59348 16192 59357 16232
rect 59299 16191 59357 16192
rect 59683 16232 59741 16233
rect 59683 16192 59692 16232
rect 59732 16192 59741 16232
rect 59683 16191 59741 16192
rect 60067 16232 60125 16233
rect 60067 16192 60076 16232
rect 60116 16192 60125 16232
rect 60067 16191 60125 16192
rect 60547 16232 60605 16233
rect 60547 16192 60556 16232
rect 60596 16192 60605 16232
rect 60547 16191 60605 16192
rect 61411 16232 61469 16233
rect 61411 16192 61420 16232
rect 61460 16192 61469 16232
rect 61411 16191 61469 16192
rect 62083 16232 62141 16233
rect 62083 16192 62092 16232
rect 62132 16192 62141 16232
rect 62083 16191 62141 16192
rect 62371 16232 62429 16233
rect 62371 16192 62380 16232
rect 62420 16192 62429 16232
rect 62371 16191 62429 16192
rect 62659 16232 62717 16233
rect 62659 16192 62668 16232
rect 62708 16192 62717 16232
rect 62659 16191 62717 16192
rect 62947 16232 63005 16233
rect 62947 16192 62956 16232
rect 62996 16192 63005 16232
rect 62947 16191 63005 16192
rect 63235 16232 63293 16233
rect 63235 16192 63244 16232
rect 63284 16192 63293 16232
rect 63235 16191 63293 16192
rect 63523 16232 63581 16233
rect 63523 16192 63532 16232
rect 63572 16192 63581 16232
rect 63523 16191 63581 16192
rect 63811 16232 63869 16233
rect 63811 16192 63820 16232
rect 63860 16192 63869 16232
rect 63811 16191 63869 16192
rect 64099 16232 64157 16233
rect 64099 16192 64108 16232
rect 64148 16192 64157 16232
rect 64099 16191 64157 16192
rect 64483 16232 64541 16233
rect 64483 16192 64492 16232
rect 64532 16192 64541 16232
rect 64483 16191 64541 16192
rect 64963 16232 65021 16233
rect 64963 16192 64972 16232
rect 65012 16192 65021 16232
rect 64963 16191 65021 16192
rect 65347 16232 65405 16233
rect 65347 16192 65356 16232
rect 65396 16192 65405 16232
rect 65347 16191 65405 16192
rect 65731 16232 65789 16233
rect 65731 16192 65740 16232
rect 65780 16192 65789 16232
rect 65731 16191 65789 16192
rect 66115 16232 66173 16233
rect 66115 16192 66124 16232
rect 66164 16192 66173 16232
rect 66115 16191 66173 16192
rect 66499 16232 66557 16233
rect 66499 16192 66508 16232
rect 66548 16192 66557 16232
rect 66499 16191 66557 16192
rect 66979 16232 67037 16233
rect 66979 16192 66988 16232
rect 67028 16192 67037 16232
rect 66979 16191 67037 16192
rect 67363 16232 67421 16233
rect 67363 16192 67372 16232
rect 67412 16192 67421 16232
rect 67363 16191 67421 16192
rect 67747 16232 67805 16233
rect 67747 16192 67756 16232
rect 67796 16192 67805 16232
rect 67747 16191 67805 16192
rect 68131 16232 68189 16233
rect 68131 16192 68140 16232
rect 68180 16192 68189 16232
rect 68131 16191 68189 16192
rect 68515 16232 68573 16233
rect 68515 16192 68524 16232
rect 68564 16192 68573 16232
rect 68515 16191 68573 16192
rect 68995 16232 69053 16233
rect 68995 16192 69004 16232
rect 69044 16192 69053 16232
rect 68995 16191 69053 16192
rect 69379 16232 69437 16233
rect 69379 16192 69388 16232
rect 69428 16192 69437 16232
rect 69379 16191 69437 16192
rect 69763 16232 69821 16233
rect 69763 16192 69772 16232
rect 69812 16192 69821 16232
rect 69763 16191 69821 16192
rect 70147 16232 70205 16233
rect 70147 16192 70156 16232
rect 70196 16192 70205 16232
rect 70915 16232 70973 16233
rect 70147 16191 70205 16192
rect 70526 16221 70568 16230
rect 53268 16170 53310 16179
rect 70526 16181 70527 16221
rect 70567 16181 70568 16221
rect 70915 16192 70924 16232
rect 70964 16192 70973 16232
rect 70915 16191 70973 16192
rect 71299 16232 71357 16233
rect 71299 16192 71308 16232
rect 71348 16192 71357 16232
rect 71299 16191 71357 16192
rect 71779 16232 71837 16233
rect 71779 16192 71788 16232
rect 71828 16192 71837 16232
rect 71779 16191 71837 16192
rect 72163 16232 72221 16233
rect 72163 16192 72172 16232
rect 72212 16192 72221 16232
rect 72163 16191 72221 16192
rect 72547 16232 72605 16233
rect 72547 16192 72556 16232
rect 72596 16192 72605 16232
rect 72547 16191 72605 16192
rect 72931 16232 72989 16233
rect 72931 16192 72940 16232
rect 72980 16192 72989 16232
rect 72931 16191 72989 16192
rect 73315 16232 73373 16233
rect 73315 16192 73324 16232
rect 73364 16192 73373 16232
rect 73315 16191 73373 16192
rect 73699 16232 73757 16233
rect 73699 16192 73708 16232
rect 73748 16192 73757 16232
rect 73699 16191 73757 16192
rect 74179 16232 74237 16233
rect 74179 16192 74188 16232
rect 74228 16192 74237 16232
rect 74179 16191 74237 16192
rect 74563 16232 74621 16233
rect 74563 16192 74572 16232
rect 74612 16192 74621 16232
rect 74563 16191 74621 16192
rect 74947 16232 75005 16233
rect 74947 16192 74956 16232
rect 74996 16192 75005 16232
rect 74947 16191 75005 16192
rect 75331 16232 75389 16233
rect 75331 16192 75340 16232
rect 75380 16192 75389 16232
rect 75331 16191 75389 16192
rect 75715 16232 75773 16233
rect 75715 16192 75724 16232
rect 75764 16192 75773 16232
rect 75715 16191 75773 16192
rect 76579 16232 76637 16233
rect 76579 16192 76588 16232
rect 76628 16192 76637 16232
rect 76579 16191 76637 16192
rect 76963 16232 77021 16233
rect 76963 16192 76972 16232
rect 77012 16192 77021 16232
rect 76963 16191 77021 16192
rect 77155 16232 77213 16233
rect 77155 16192 77164 16232
rect 77204 16192 77213 16232
rect 77155 16191 77213 16192
rect 77443 16232 77501 16233
rect 77443 16192 77452 16232
rect 77492 16192 77501 16232
rect 77443 16191 77501 16192
rect 77827 16232 77885 16233
rect 77827 16192 77836 16232
rect 77876 16192 77885 16232
rect 77827 16191 77885 16192
rect 78211 16232 78269 16233
rect 78211 16192 78220 16232
rect 78260 16192 78269 16232
rect 78211 16191 78269 16192
rect 78595 16232 78653 16233
rect 78595 16192 78604 16232
rect 78644 16192 78653 16232
rect 78595 16191 78653 16192
rect 78883 16232 78941 16233
rect 78883 16192 78892 16232
rect 78932 16192 78941 16232
rect 78883 16191 78941 16192
rect 79171 16232 79229 16233
rect 79171 16192 79180 16232
rect 79220 16192 79229 16232
rect 79171 16191 79229 16192
rect 70526 16172 70568 16181
rect 3435 16148 3477 16157
rect 3435 16108 3436 16148
rect 3476 16108 3477 16148
rect 3435 16099 3477 16108
rect 4587 16148 4629 16157
rect 4587 16108 4588 16148
rect 4628 16108 4629 16148
rect 4587 16099 4629 16108
rect 27435 16148 27477 16157
rect 27435 16108 27436 16148
rect 27476 16108 27477 16148
rect 27435 16099 27477 16108
rect 30987 16148 31029 16157
rect 30987 16108 30988 16148
rect 31028 16108 31029 16148
rect 30987 16099 31029 16108
rect 34059 16148 34101 16157
rect 34059 16108 34060 16148
rect 34100 16108 34101 16148
rect 34059 16099 34101 16108
rect 37035 16148 37077 16157
rect 37035 16108 37036 16148
rect 37076 16108 37077 16148
rect 37035 16099 37077 16108
rect 40011 16148 40053 16157
rect 40011 16108 40012 16148
rect 40052 16108 40053 16148
rect 40011 16099 40053 16108
rect 40299 16148 40341 16157
rect 40299 16108 40300 16148
rect 40340 16108 40341 16148
rect 40299 16099 40341 16108
rect 43275 16148 43317 16157
rect 43275 16108 43276 16148
rect 43316 16108 43317 16148
rect 43275 16099 43317 16108
rect 55371 16148 55413 16157
rect 55371 16108 55372 16148
rect 55412 16108 55413 16148
rect 55371 16099 55413 16108
rect 2187 16064 2229 16073
rect 2187 16024 2188 16064
rect 2228 16024 2229 16064
rect 2187 16015 2229 16024
rect 2955 16064 2997 16073
rect 2955 16024 2956 16064
rect 2996 16024 2997 16064
rect 2955 16015 2997 16024
rect 6979 16064 7037 16065
rect 6979 16024 6988 16064
rect 7028 16024 7037 16064
rect 6979 16023 7037 16024
rect 33379 16064 33437 16065
rect 33379 16024 33388 16064
rect 33428 16024 33437 16064
rect 33379 16023 33437 16024
rect 45667 16064 45725 16065
rect 45667 16024 45676 16064
rect 45716 16024 45725 16064
rect 45667 16023 45725 16024
rect 46443 16064 46485 16073
rect 46443 16024 46444 16064
rect 46484 16024 46485 16064
rect 46443 16015 46485 16024
rect 51043 16064 51101 16065
rect 51043 16024 51052 16064
rect 51092 16024 51101 16064
rect 51043 16023 51101 16024
rect 52675 16064 52733 16065
rect 52675 16024 52684 16064
rect 52724 16024 52733 16064
rect 52675 16023 52733 16024
rect 57003 16064 57045 16073
rect 57003 16024 57004 16064
rect 57044 16024 57045 16064
rect 57003 16015 57045 16024
rect 59019 16064 59061 16073
rect 59019 16024 59020 16064
rect 59060 16024 59061 16064
rect 59019 16015 59061 16024
rect 59403 16064 59445 16073
rect 59403 16024 59404 16064
rect 59444 16024 59445 16064
rect 59403 16015 59445 16024
rect 59787 16064 59829 16073
rect 59787 16024 59788 16064
rect 59828 16024 59829 16064
rect 59787 16015 59829 16024
rect 61899 16064 61941 16073
rect 61899 16024 61900 16064
rect 61940 16024 61941 16064
rect 61899 16015 61941 16024
rect 62763 16064 62805 16073
rect 62763 16024 62764 16064
rect 62804 16024 62805 16064
rect 62763 16015 62805 16024
rect 64203 16064 64245 16073
rect 64203 16024 64204 16064
rect 64244 16024 64245 16064
rect 64203 16015 64245 16024
rect 66219 16064 66261 16073
rect 66219 16024 66220 16064
rect 66260 16024 66261 16064
rect 66219 16015 66261 16024
rect 68619 16064 68661 16073
rect 68619 16024 68620 16064
rect 68660 16024 68661 16064
rect 68619 16015 68661 16024
rect 73803 16064 73845 16073
rect 73803 16024 73804 16064
rect 73844 16024 73845 16064
rect 73803 16015 73845 16024
rect 576 15896 79584 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 79584 15896
rect 576 15832 79584 15856
rect 3627 15728 3669 15737
rect 3627 15688 3628 15728
rect 3668 15688 3669 15728
rect 3627 15679 3669 15688
rect 4387 15728 4445 15729
rect 4387 15688 4396 15728
rect 4436 15688 4445 15728
rect 4387 15687 4445 15688
rect 33859 15728 33917 15729
rect 33859 15688 33868 15728
rect 33908 15688 33917 15728
rect 33859 15687 33917 15688
rect 34915 15728 34973 15729
rect 34915 15688 34924 15728
rect 34964 15688 34973 15728
rect 34915 15687 34973 15688
rect 40483 15728 40541 15729
rect 40483 15688 40492 15728
rect 40532 15688 40541 15728
rect 40483 15687 40541 15688
rect 45955 15728 46013 15729
rect 45955 15688 45964 15728
rect 46004 15688 46013 15728
rect 45955 15687 46013 15688
rect 49699 15728 49757 15729
rect 49699 15688 49708 15728
rect 49748 15688 49757 15728
rect 49699 15687 49757 15688
rect 59491 15728 59549 15729
rect 59491 15688 59500 15728
rect 59540 15688 59549 15728
rect 59491 15687 59549 15688
rect 67843 15728 67901 15729
rect 67843 15688 67852 15728
rect 67892 15688 67901 15728
rect 67843 15687 67901 15688
rect 70539 15728 70581 15737
rect 70539 15688 70540 15728
rect 70580 15688 70581 15728
rect 70539 15679 70581 15688
rect 79467 15728 79509 15737
rect 79467 15688 79468 15728
rect 79508 15688 79509 15728
rect 79467 15679 79509 15688
rect 53163 15644 53205 15653
rect 53163 15604 53164 15644
rect 53204 15604 53205 15644
rect 53163 15595 53205 15604
rect 1035 15560 1077 15569
rect 1035 15520 1036 15560
rect 1076 15520 1077 15560
rect 1035 15511 1077 15520
rect 1411 15560 1469 15561
rect 1411 15520 1420 15560
rect 1460 15520 1469 15560
rect 1411 15519 1469 15520
rect 2275 15560 2333 15561
rect 2275 15520 2284 15560
rect 2324 15520 2333 15560
rect 2275 15519 2333 15520
rect 4195 15560 4253 15561
rect 4195 15520 4204 15560
rect 4244 15520 4253 15560
rect 4195 15519 4253 15520
rect 4299 15560 4341 15569
rect 4299 15520 4300 15560
rect 4340 15520 4341 15560
rect 4299 15511 4341 15520
rect 4491 15560 4533 15569
rect 4491 15520 4492 15560
rect 4532 15520 4533 15560
rect 4491 15511 4533 15520
rect 4675 15560 4733 15561
rect 4675 15520 4684 15560
rect 4724 15520 4733 15560
rect 4675 15519 4733 15520
rect 4779 15560 4821 15569
rect 4779 15520 4780 15560
rect 4820 15520 4821 15560
rect 4779 15511 4821 15520
rect 4875 15560 4917 15569
rect 4875 15520 4876 15560
rect 4916 15520 4917 15560
rect 4875 15511 4917 15520
rect 31939 15560 31997 15561
rect 31939 15520 31948 15560
rect 31988 15520 31997 15560
rect 31939 15519 31997 15520
rect 32139 15560 32181 15569
rect 32139 15520 32140 15560
rect 32180 15520 32181 15560
rect 32139 15511 32181 15520
rect 32811 15560 32853 15569
rect 32811 15520 32812 15560
rect 32852 15520 32853 15560
rect 32811 15511 32853 15520
rect 33003 15560 33045 15569
rect 33003 15520 33004 15560
rect 33044 15520 33045 15560
rect 33003 15511 33045 15520
rect 33117 15560 33159 15569
rect 33117 15520 33118 15560
rect 33158 15520 33159 15560
rect 33117 15511 33159 15520
rect 33291 15560 33333 15569
rect 33291 15520 33292 15560
rect 33332 15520 33333 15560
rect 33291 15511 33333 15520
rect 33387 15560 33429 15569
rect 33387 15520 33388 15560
rect 33428 15520 33429 15560
rect 33387 15511 33429 15520
rect 33483 15560 33525 15569
rect 33483 15520 33484 15560
rect 33524 15520 33525 15560
rect 33483 15511 33525 15520
rect 33579 15560 33621 15569
rect 33579 15520 33580 15560
rect 33620 15520 33621 15560
rect 33579 15511 33621 15520
rect 33771 15560 33813 15569
rect 33771 15520 33772 15560
rect 33812 15520 33813 15560
rect 33771 15511 33813 15520
rect 33963 15560 34005 15569
rect 33963 15520 33964 15560
rect 34004 15520 34005 15560
rect 33963 15511 34005 15520
rect 34051 15560 34109 15561
rect 34051 15520 34060 15560
rect 34100 15520 34109 15560
rect 34051 15519 34109 15520
rect 34443 15560 34485 15569
rect 34443 15520 34444 15560
rect 34484 15520 34485 15560
rect 34443 15511 34485 15520
rect 34635 15560 34677 15569
rect 34635 15520 34636 15560
rect 34676 15520 34677 15560
rect 34635 15511 34677 15520
rect 34723 15560 34781 15561
rect 34723 15520 34732 15560
rect 34772 15520 34781 15560
rect 34723 15519 34781 15520
rect 36067 15560 36125 15561
rect 36067 15520 36076 15560
rect 36116 15520 36125 15560
rect 36067 15519 36125 15520
rect 36931 15560 36989 15561
rect 36931 15520 36940 15560
rect 36980 15520 36989 15560
rect 36931 15519 36989 15520
rect 37323 15560 37365 15569
rect 37323 15520 37324 15560
rect 37364 15520 37365 15560
rect 37323 15511 37365 15520
rect 37515 15560 37557 15569
rect 37515 15520 37516 15560
rect 37556 15520 37557 15560
rect 37515 15511 37557 15520
rect 37707 15560 37749 15569
rect 37707 15520 37708 15560
rect 37748 15520 37749 15560
rect 37707 15511 37749 15520
rect 37795 15560 37853 15561
rect 37795 15520 37804 15560
rect 37844 15520 37853 15560
rect 37795 15519 37853 15520
rect 39051 15560 39093 15569
rect 39051 15520 39052 15560
rect 39092 15520 39093 15560
rect 39051 15511 39093 15520
rect 39147 15560 39189 15569
rect 39147 15520 39148 15560
rect 39188 15520 39189 15560
rect 39147 15511 39189 15520
rect 39235 15560 39293 15561
rect 39235 15520 39244 15560
rect 39284 15520 39293 15560
rect 39235 15519 39293 15520
rect 39723 15560 39765 15569
rect 39723 15520 39724 15560
rect 39764 15520 39765 15560
rect 39723 15511 39765 15520
rect 39819 15560 39861 15569
rect 39819 15520 39820 15560
rect 39860 15520 39861 15560
rect 39819 15511 39861 15520
rect 40099 15560 40157 15561
rect 40099 15520 40108 15560
rect 40148 15520 40157 15560
rect 40099 15519 40157 15520
rect 40395 15560 40437 15569
rect 40395 15520 40396 15560
rect 40436 15520 40437 15560
rect 40395 15511 40437 15520
rect 40587 15560 40629 15569
rect 40587 15520 40588 15560
rect 40628 15520 40629 15560
rect 40587 15511 40629 15520
rect 40675 15560 40733 15561
rect 40675 15520 40684 15560
rect 40724 15520 40733 15560
rect 40675 15519 40733 15520
rect 41835 15560 41877 15569
rect 41835 15520 41836 15560
rect 41876 15520 41877 15560
rect 41835 15511 41877 15520
rect 42027 15560 42069 15569
rect 42027 15520 42028 15560
rect 42068 15520 42069 15560
rect 42027 15511 42069 15520
rect 42115 15560 42173 15561
rect 42115 15520 42124 15560
rect 42164 15520 42173 15560
rect 42115 15519 42173 15520
rect 45387 15560 45429 15569
rect 45387 15520 45388 15560
rect 45428 15520 45429 15560
rect 45387 15511 45429 15520
rect 45483 15560 45525 15569
rect 45483 15520 45484 15560
rect 45524 15520 45525 15560
rect 45483 15511 45525 15520
rect 45579 15560 45621 15569
rect 45579 15520 45580 15560
rect 45620 15520 45621 15560
rect 45579 15511 45621 15520
rect 45675 15560 45717 15569
rect 45675 15520 45676 15560
rect 45716 15520 45717 15560
rect 45675 15511 45717 15520
rect 45867 15560 45909 15569
rect 45867 15520 45868 15560
rect 45908 15520 45909 15560
rect 45867 15511 45909 15520
rect 46059 15560 46101 15569
rect 46059 15520 46060 15560
rect 46100 15520 46101 15560
rect 46059 15511 46101 15520
rect 46147 15560 46205 15561
rect 46147 15520 46156 15560
rect 46196 15520 46205 15560
rect 46147 15519 46205 15520
rect 46347 15560 46389 15569
rect 46347 15520 46348 15560
rect 46388 15520 46389 15560
rect 46347 15511 46389 15520
rect 46443 15560 46485 15569
rect 46443 15520 46444 15560
rect 46484 15520 46485 15560
rect 46443 15511 46485 15520
rect 46531 15560 46589 15561
rect 46531 15520 46540 15560
rect 46580 15520 46589 15560
rect 46531 15519 46589 15520
rect 46915 15560 46973 15561
rect 46915 15520 46924 15560
rect 46964 15520 46973 15560
rect 47307 15560 47349 15569
rect 46915 15519 46973 15520
rect 47211 15518 47253 15527
rect 47211 15478 47212 15518
rect 47252 15478 47253 15518
rect 47307 15520 47308 15560
rect 47348 15520 47349 15560
rect 47307 15511 47349 15520
rect 47787 15560 47829 15569
rect 47787 15520 47788 15560
rect 47828 15520 47829 15560
rect 47787 15511 47829 15520
rect 47971 15560 48029 15561
rect 47971 15520 47980 15560
rect 48020 15520 48029 15560
rect 47971 15519 48029 15520
rect 49803 15560 49845 15569
rect 49803 15520 49804 15560
rect 49844 15520 49845 15560
rect 49803 15511 49845 15520
rect 49899 15560 49941 15569
rect 49899 15520 49900 15560
rect 49940 15520 49941 15560
rect 49899 15511 49941 15520
rect 49995 15560 50037 15569
rect 49995 15520 49996 15560
rect 50036 15520 50037 15560
rect 50841 15567 50899 15568
rect 50841 15527 50850 15567
rect 50890 15527 50899 15567
rect 50841 15526 50899 15527
rect 50955 15560 50997 15569
rect 49995 15511 50037 15520
rect 50955 15520 50956 15560
rect 50996 15520 50997 15560
rect 50955 15511 50997 15520
rect 51147 15560 51189 15569
rect 51147 15520 51148 15560
rect 51188 15520 51189 15560
rect 51147 15511 51189 15520
rect 51531 15560 51573 15569
rect 51531 15520 51532 15560
rect 51572 15520 51573 15560
rect 51531 15511 51573 15520
rect 51627 15560 51669 15569
rect 51627 15520 51628 15560
rect 51668 15520 51669 15560
rect 51627 15511 51669 15520
rect 51723 15560 51765 15569
rect 51723 15520 51724 15560
rect 51764 15520 51765 15560
rect 51723 15511 51765 15520
rect 51819 15560 51861 15569
rect 51819 15520 51820 15560
rect 51860 15520 51861 15560
rect 51819 15511 51861 15520
rect 52195 15560 52253 15561
rect 52195 15520 52204 15560
rect 52244 15520 52253 15560
rect 52195 15519 52253 15520
rect 52491 15560 52533 15569
rect 52491 15520 52492 15560
rect 52532 15520 52533 15560
rect 52491 15511 52533 15520
rect 52587 15560 52629 15569
rect 52587 15520 52588 15560
rect 52628 15520 52629 15560
rect 52587 15511 52629 15520
rect 53539 15560 53597 15561
rect 53539 15520 53548 15560
rect 53588 15520 53597 15560
rect 53539 15519 53597 15520
rect 54403 15560 54461 15561
rect 54403 15520 54412 15560
rect 54452 15520 54461 15560
rect 54403 15519 54461 15520
rect 57099 15560 57141 15569
rect 57099 15520 57100 15560
rect 57140 15520 57141 15560
rect 57099 15511 57141 15520
rect 57475 15560 57533 15561
rect 57475 15520 57484 15560
rect 57524 15520 57533 15560
rect 57475 15519 57533 15520
rect 58339 15560 58397 15561
rect 58339 15520 58348 15560
rect 58388 15520 58397 15560
rect 58339 15519 58397 15520
rect 60555 15560 60597 15569
rect 60555 15520 60556 15560
rect 60596 15520 60597 15560
rect 60555 15511 60597 15520
rect 60931 15560 60989 15561
rect 60931 15520 60940 15560
rect 60980 15520 60989 15560
rect 60931 15519 60989 15520
rect 61795 15560 61853 15561
rect 61795 15520 61804 15560
rect 61844 15520 61853 15560
rect 61795 15519 61853 15520
rect 64779 15560 64821 15569
rect 64779 15520 64780 15560
rect 64820 15520 64821 15560
rect 64779 15511 64821 15520
rect 64963 15560 65021 15561
rect 64963 15520 64972 15560
rect 65012 15520 65021 15560
rect 64963 15519 65021 15520
rect 65451 15560 65493 15569
rect 65451 15520 65452 15560
rect 65492 15520 65493 15560
rect 65451 15511 65493 15520
rect 65827 15560 65885 15561
rect 65827 15520 65836 15560
rect 65876 15520 65885 15560
rect 65827 15519 65885 15520
rect 66691 15560 66749 15561
rect 66691 15520 66700 15560
rect 66740 15520 66749 15560
rect 66691 15519 66749 15520
rect 70051 15560 70109 15561
rect 70051 15520 70060 15560
rect 70100 15520 70109 15560
rect 70051 15519 70109 15520
rect 70155 15560 70197 15569
rect 70155 15520 70156 15560
rect 70196 15520 70197 15560
rect 70155 15511 70197 15520
rect 70347 15560 70389 15569
rect 70347 15520 70348 15560
rect 70388 15520 70389 15560
rect 70347 15511 70389 15520
rect 75139 15560 75197 15561
rect 75139 15520 75148 15560
rect 75188 15520 75197 15560
rect 75139 15519 75197 15520
rect 75339 15560 75381 15569
rect 75339 15520 75340 15560
rect 75380 15520 75381 15560
rect 75339 15511 75381 15520
rect 79363 15560 79421 15561
rect 79363 15520 79372 15560
rect 79412 15520 79421 15560
rect 79363 15519 79421 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 3811 15476 3869 15477
rect 3811 15436 3820 15476
rect 3860 15436 3869 15476
rect 47211 15469 47253 15478
rect 55563 15476 55605 15485
rect 3811 15435 3869 15436
rect 55563 15436 55564 15476
rect 55604 15436 55605 15476
rect 55563 15427 55605 15436
rect 68707 15476 68765 15477
rect 68707 15436 68716 15476
rect 68756 15436 68765 15476
rect 68707 15435 68765 15436
rect 69859 15476 69917 15477
rect 69859 15436 69868 15476
rect 69908 15436 69917 15476
rect 69859 15435 69917 15436
rect 70723 15476 70781 15477
rect 70723 15436 70732 15476
rect 70772 15436 70781 15476
rect 70723 15435 70781 15436
rect 71107 15476 71165 15477
rect 71107 15436 71116 15476
rect 71156 15436 71165 15476
rect 71107 15435 71165 15436
rect 5067 15392 5109 15401
rect 5067 15352 5068 15392
rect 5108 15352 5109 15392
rect 5067 15343 5109 15352
rect 31467 15392 31509 15401
rect 31467 15352 31468 15392
rect 31508 15352 31509 15392
rect 31467 15343 31509 15352
rect 34443 15392 34485 15401
rect 34443 15352 34444 15392
rect 34484 15352 34485 15392
rect 34443 15343 34485 15352
rect 37515 15392 37557 15401
rect 37515 15352 37516 15392
rect 37556 15352 37557 15392
rect 37515 15343 37557 15352
rect 38187 15392 38229 15401
rect 38187 15352 38188 15392
rect 38228 15352 38229 15392
rect 38187 15343 38229 15352
rect 39427 15392 39485 15393
rect 39427 15352 39436 15392
rect 39476 15352 39485 15392
rect 39427 15351 39485 15352
rect 40875 15392 40917 15401
rect 40875 15352 40876 15392
rect 40916 15352 40917 15392
rect 40875 15343 40917 15352
rect 43755 15392 43797 15401
rect 43755 15352 43756 15392
rect 43796 15352 43797 15392
rect 43755 15343 43797 15352
rect 48459 15392 48501 15401
rect 48459 15352 48460 15392
rect 48500 15352 48501 15392
rect 48459 15343 48501 15352
rect 49131 15392 49173 15401
rect 49131 15352 49132 15392
rect 49172 15352 49173 15392
rect 49131 15343 49173 15352
rect 68043 15392 68085 15401
rect 68043 15352 68044 15392
rect 68084 15352 68085 15392
rect 68043 15343 68085 15352
rect 71307 15392 71349 15401
rect 71307 15352 71308 15392
rect 71348 15352 71349 15392
rect 71307 15343 71349 15352
rect 72651 15392 72693 15401
rect 72651 15352 72652 15392
rect 72692 15352 72693 15392
rect 72651 15343 72693 15352
rect 76683 15392 76725 15401
rect 76683 15352 76684 15392
rect 76724 15352 76725 15392
rect 76683 15343 76725 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 3427 15308 3485 15309
rect 3427 15268 3436 15308
rect 3476 15268 3485 15308
rect 3427 15267 3485 15268
rect 3627 15308 3669 15317
rect 3627 15268 3628 15308
rect 3668 15268 3669 15308
rect 3627 15259 3669 15268
rect 32043 15308 32085 15317
rect 32043 15268 32044 15308
rect 32084 15268 32085 15308
rect 32043 15259 32085 15268
rect 32811 15308 32853 15317
rect 32811 15268 32812 15308
rect 32852 15268 32853 15308
rect 32811 15259 32853 15268
rect 41835 15308 41877 15317
rect 41835 15268 41836 15308
rect 41876 15268 41877 15308
rect 41835 15259 41877 15268
rect 47587 15308 47645 15309
rect 47587 15268 47596 15308
rect 47636 15268 47645 15308
rect 47587 15267 47645 15268
rect 47883 15308 47925 15317
rect 47883 15268 47884 15308
rect 47924 15268 47925 15308
rect 47883 15259 47925 15268
rect 51147 15308 51189 15317
rect 51147 15268 51148 15308
rect 51188 15268 51189 15308
rect 51147 15259 51189 15268
rect 52867 15308 52925 15309
rect 52867 15268 52876 15308
rect 52916 15268 52925 15308
rect 52867 15267 52925 15268
rect 59491 15308 59549 15309
rect 59491 15268 59500 15308
rect 59540 15268 59549 15308
rect 59491 15267 59549 15268
rect 62947 15308 63005 15309
rect 62947 15268 62956 15308
rect 62996 15268 63005 15308
rect 62947 15267 63005 15268
rect 64875 15308 64917 15317
rect 64875 15268 64876 15308
rect 64916 15268 64917 15308
rect 64875 15259 64917 15268
rect 68907 15308 68949 15317
rect 68907 15268 68908 15308
rect 68948 15268 68949 15308
rect 68907 15259 68949 15268
rect 69675 15308 69717 15317
rect 69675 15268 69676 15308
rect 69716 15268 69717 15308
rect 69675 15259 69717 15268
rect 70347 15308 70389 15317
rect 70347 15268 70348 15308
rect 70388 15268 70389 15308
rect 70347 15259 70389 15268
rect 70923 15308 70965 15317
rect 70923 15268 70924 15308
rect 70964 15268 70965 15308
rect 70923 15259 70965 15268
rect 75243 15308 75285 15317
rect 75243 15268 75244 15308
rect 75284 15268 75285 15308
rect 75243 15259 75285 15268
rect 576 15140 79584 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 75112 15140
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75480 15100 79584 15140
rect 576 15076 79584 15100
rect 1995 14972 2037 14981
rect 1995 14932 1996 14972
rect 2036 14932 2037 14972
rect 1995 14923 2037 14932
rect 3235 14972 3293 14973
rect 3235 14932 3244 14972
rect 3284 14932 3293 14972
rect 3235 14931 3293 14932
rect 45579 14972 45621 14981
rect 45579 14932 45580 14972
rect 45620 14932 45621 14972
rect 45579 14923 45621 14932
rect 50371 14972 50429 14973
rect 50371 14932 50380 14972
rect 50420 14932 50429 14972
rect 50371 14931 50429 14932
rect 53155 14972 53213 14973
rect 53155 14932 53164 14972
rect 53204 14932 53213 14972
rect 53155 14931 53213 14932
rect 56907 14972 56949 14981
rect 56907 14932 56908 14972
rect 56948 14932 56949 14972
rect 56907 14923 56949 14932
rect 60939 14972 60981 14981
rect 60939 14932 60940 14972
rect 60980 14932 60981 14972
rect 60939 14923 60981 14932
rect 65355 14972 65397 14981
rect 65355 14932 65356 14972
rect 65396 14932 65397 14972
rect 65355 14923 65397 14932
rect 72739 14972 72797 14973
rect 72739 14932 72748 14972
rect 72788 14932 72797 14972
rect 72739 14931 72797 14932
rect 75331 14972 75389 14973
rect 75331 14932 75340 14972
rect 75380 14932 75389 14972
rect 75331 14931 75389 14932
rect 78595 14972 78653 14973
rect 78595 14932 78604 14972
rect 78644 14932 78653 14972
rect 78595 14931 78653 14932
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 33483 14888 33525 14897
rect 33483 14848 33484 14888
rect 33524 14848 33525 14888
rect 33483 14839 33525 14848
rect 35595 14888 35637 14897
rect 35595 14848 35596 14888
rect 35636 14848 35637 14888
rect 35595 14839 35637 14848
rect 40011 14888 40053 14897
rect 40011 14848 40012 14888
rect 40052 14848 40053 14888
rect 40011 14839 40053 14848
rect 45099 14888 45141 14897
rect 45099 14848 45100 14888
rect 45140 14848 45141 14888
rect 45099 14839 45141 14848
rect 54315 14888 54357 14897
rect 54315 14848 54316 14888
rect 54356 14848 54357 14888
rect 54315 14839 54357 14848
rect 56707 14888 56765 14889
rect 56707 14848 56716 14888
rect 56756 14848 56765 14888
rect 56707 14847 56765 14848
rect 57483 14888 57525 14897
rect 57483 14848 57484 14888
rect 57524 14848 57525 14888
rect 57483 14839 57525 14848
rect 58635 14888 58677 14897
rect 58635 14848 58636 14888
rect 58676 14848 58677 14888
rect 58635 14839 58677 14848
rect 61419 14888 61461 14897
rect 61419 14848 61420 14888
rect 61460 14848 61461 14888
rect 61419 14839 61461 14848
rect 64099 14888 64157 14889
rect 64099 14848 64108 14888
rect 64148 14848 64157 14888
rect 64099 14847 64157 14848
rect 65931 14888 65973 14897
rect 65931 14848 65932 14888
rect 65972 14848 65973 14888
rect 65931 14839 65973 14848
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 1219 14804 1277 14805
rect 1219 14764 1228 14804
rect 1268 14764 1277 14804
rect 60739 14804 60797 14805
rect 1219 14763 1277 14764
rect 2859 14762 2901 14771
rect 60739 14764 60748 14804
rect 60788 14764 60797 14804
rect 60739 14763 60797 14764
rect 61603 14804 61661 14805
rect 61603 14764 61612 14804
rect 61652 14764 61661 14804
rect 61603 14763 61661 14764
rect 61987 14804 62045 14805
rect 61987 14764 61996 14804
rect 62036 14764 62045 14804
rect 61987 14763 62045 14764
rect 62755 14804 62813 14805
rect 62755 14764 62764 14804
rect 62804 14764 62813 14804
rect 62755 14763 62813 14764
rect 67171 14804 67229 14805
rect 67171 14764 67180 14804
rect 67220 14764 67229 14804
rect 67171 14763 67229 14764
rect 1515 14720 1557 14729
rect 1515 14680 1516 14720
rect 1556 14680 1557 14720
rect 1515 14671 1557 14680
rect 1611 14720 1653 14729
rect 1611 14680 1612 14720
rect 1652 14680 1653 14720
rect 1611 14671 1653 14680
rect 1707 14720 1749 14729
rect 1707 14680 1708 14720
rect 1748 14680 1749 14720
rect 1707 14671 1749 14680
rect 1803 14720 1845 14729
rect 1803 14680 1804 14720
rect 1844 14680 1845 14720
rect 1803 14671 1845 14680
rect 1995 14720 2037 14729
rect 1995 14680 1996 14720
rect 2036 14680 2037 14720
rect 1995 14671 2037 14680
rect 2187 14720 2229 14729
rect 2859 14722 2860 14762
rect 2900 14722 2901 14762
rect 2187 14680 2188 14720
rect 2228 14680 2229 14720
rect 2187 14671 2229 14680
rect 2275 14720 2333 14721
rect 2275 14680 2284 14720
rect 2324 14680 2333 14720
rect 2275 14679 2333 14680
rect 2563 14720 2621 14721
rect 2563 14680 2572 14720
rect 2612 14680 2621 14720
rect 2859 14713 2901 14722
rect 2955 14720 2997 14729
rect 2563 14679 2621 14680
rect 2955 14680 2956 14720
rect 2996 14680 2997 14720
rect 2955 14671 2997 14680
rect 5059 14720 5117 14721
rect 5059 14680 5068 14720
rect 5108 14680 5117 14720
rect 5059 14679 5117 14680
rect 5259 14720 5301 14729
rect 5259 14680 5260 14720
rect 5300 14680 5301 14720
rect 5259 14671 5301 14680
rect 30307 14720 30365 14721
rect 30307 14680 30316 14720
rect 30356 14680 30365 14720
rect 30307 14679 30365 14680
rect 31171 14720 31229 14721
rect 31171 14680 31180 14720
rect 31220 14680 31229 14720
rect 31171 14679 31229 14680
rect 32811 14720 32853 14729
rect 32811 14680 32812 14720
rect 32852 14680 32853 14720
rect 32811 14671 32853 14680
rect 32907 14720 32949 14729
rect 32907 14680 32908 14720
rect 32948 14680 32949 14720
rect 35979 14720 36021 14729
rect 32907 14671 32949 14680
rect 33003 14699 33045 14708
rect 33003 14659 33004 14699
rect 33044 14659 33045 14699
rect 35979 14680 35980 14720
rect 36020 14680 36021 14720
rect 35979 14671 36021 14680
rect 36075 14720 36117 14729
rect 36075 14680 36076 14720
rect 36116 14680 36117 14720
rect 36075 14671 36117 14680
rect 36171 14720 36213 14729
rect 36171 14680 36172 14720
rect 36212 14680 36213 14720
rect 36171 14671 36213 14680
rect 36267 14720 36309 14729
rect 36267 14680 36268 14720
rect 36308 14680 36309 14720
rect 36267 14671 36309 14680
rect 36843 14720 36885 14729
rect 36843 14680 36844 14720
rect 36884 14680 36885 14720
rect 36843 14671 36885 14680
rect 38563 14720 38621 14721
rect 38563 14680 38572 14720
rect 38612 14680 38621 14720
rect 38563 14679 38621 14680
rect 39427 14720 39485 14721
rect 39427 14680 39436 14720
rect 39476 14680 39485 14720
rect 39427 14679 39485 14680
rect 39819 14720 39861 14729
rect 39819 14680 39820 14720
rect 39860 14680 39861 14720
rect 39819 14671 39861 14680
rect 40011 14720 40053 14729
rect 40011 14680 40012 14720
rect 40052 14680 40053 14720
rect 40011 14671 40053 14680
rect 40203 14720 40245 14729
rect 40203 14680 40204 14720
rect 40244 14680 40245 14720
rect 40203 14671 40245 14680
rect 40291 14720 40349 14721
rect 40291 14680 40300 14720
rect 40340 14680 40349 14720
rect 40291 14679 40349 14680
rect 41259 14720 41301 14729
rect 41259 14680 41260 14720
rect 41300 14680 41301 14720
rect 41259 14671 41301 14680
rect 41355 14720 41397 14729
rect 41355 14680 41356 14720
rect 41396 14680 41397 14720
rect 41355 14671 41397 14680
rect 41451 14720 41493 14729
rect 41451 14680 41452 14720
rect 41492 14680 41493 14720
rect 41451 14671 41493 14680
rect 42795 14720 42837 14729
rect 42795 14680 42796 14720
rect 42836 14680 42837 14720
rect 42795 14671 42837 14680
rect 42987 14720 43029 14729
rect 42987 14680 42988 14720
rect 43028 14680 43029 14720
rect 42987 14671 43029 14680
rect 43075 14720 43133 14721
rect 43075 14680 43084 14720
rect 43124 14680 43133 14720
rect 43075 14679 43133 14680
rect 43267 14720 43325 14721
rect 43267 14680 43276 14720
rect 43316 14680 43325 14720
rect 43267 14679 43325 14680
rect 43371 14720 43413 14729
rect 43371 14680 43372 14720
rect 43412 14680 43413 14720
rect 43371 14671 43413 14680
rect 43467 14720 43509 14729
rect 43467 14680 43468 14720
rect 43508 14680 43509 14720
rect 43467 14671 43509 14680
rect 45579 14720 45621 14729
rect 45579 14680 45580 14720
rect 45620 14680 45621 14720
rect 45579 14671 45621 14680
rect 45771 14720 45813 14729
rect 45771 14680 45772 14720
rect 45812 14680 45813 14720
rect 45771 14671 45813 14680
rect 45859 14720 45917 14721
rect 45859 14680 45868 14720
rect 45908 14680 45917 14720
rect 45859 14679 45917 14680
rect 46251 14720 46293 14729
rect 46251 14680 46252 14720
rect 46292 14680 46293 14720
rect 46251 14671 46293 14680
rect 47395 14720 47453 14721
rect 47395 14680 47404 14720
rect 47444 14680 47453 14720
rect 47395 14679 47453 14680
rect 47595 14720 47637 14729
rect 47595 14680 47596 14720
rect 47636 14680 47637 14720
rect 47595 14671 47637 14680
rect 48355 14720 48413 14721
rect 48355 14680 48364 14720
rect 48404 14680 48413 14720
rect 48355 14679 48413 14680
rect 49219 14720 49277 14721
rect 49219 14680 49228 14720
rect 49268 14680 49277 14720
rect 49219 14679 49277 14680
rect 51139 14720 51197 14721
rect 51139 14680 51148 14720
rect 51188 14680 51197 14720
rect 51139 14679 51197 14680
rect 52003 14720 52061 14721
rect 52003 14680 52012 14720
rect 52052 14680 52061 14720
rect 52003 14679 52061 14680
rect 56035 14720 56093 14721
rect 56035 14680 56044 14720
rect 56084 14680 56093 14720
rect 56035 14679 56093 14680
rect 56331 14720 56373 14729
rect 56331 14680 56332 14720
rect 56372 14680 56373 14720
rect 56331 14671 56373 14680
rect 56907 14720 56949 14729
rect 56907 14680 56908 14720
rect 56948 14680 56949 14720
rect 56907 14671 56949 14680
rect 57099 14720 57141 14729
rect 57099 14680 57100 14720
rect 57140 14680 57141 14720
rect 57099 14671 57141 14680
rect 57187 14720 57245 14721
rect 57187 14680 57196 14720
rect 57236 14680 57245 14720
rect 57187 14679 57245 14680
rect 57379 14720 57437 14721
rect 57379 14680 57388 14720
rect 57428 14680 57437 14720
rect 57379 14679 57437 14680
rect 57579 14720 57621 14729
rect 57579 14680 57580 14720
rect 57620 14680 57621 14720
rect 57579 14671 57621 14680
rect 60939 14720 60981 14729
rect 60939 14680 60940 14720
rect 60980 14680 60981 14720
rect 60939 14671 60981 14680
rect 61131 14720 61173 14729
rect 61131 14680 61132 14720
rect 61172 14680 61173 14720
rect 61131 14671 61173 14680
rect 61219 14720 61277 14721
rect 61219 14680 61228 14720
rect 61268 14680 61277 14720
rect 61219 14679 61277 14680
rect 62179 14720 62237 14721
rect 62179 14680 62188 14720
rect 62228 14680 62237 14720
rect 62179 14679 62237 14680
rect 62283 14720 62325 14729
rect 62283 14680 62284 14720
rect 62324 14680 62325 14720
rect 62283 14671 62325 14680
rect 62379 14720 62421 14729
rect 62379 14680 62380 14720
rect 62420 14680 62421 14720
rect 62379 14671 62421 14680
rect 63715 14720 63773 14721
rect 63715 14680 63724 14720
rect 63764 14680 63773 14720
rect 63715 14679 63773 14680
rect 63819 14720 63861 14729
rect 63819 14680 63820 14720
rect 63860 14680 63861 14720
rect 63819 14671 63861 14680
rect 63915 14720 63957 14729
rect 63915 14680 63916 14720
rect 63956 14680 63957 14720
rect 63915 14671 63957 14680
rect 64491 14720 64533 14729
rect 64491 14680 64492 14720
rect 64532 14680 64533 14720
rect 64491 14671 64533 14680
rect 64771 14720 64829 14721
rect 64771 14680 64780 14720
rect 64820 14680 64829 14720
rect 64771 14679 64829 14680
rect 65059 14720 65117 14721
rect 65059 14680 65068 14720
rect 65108 14680 65117 14720
rect 65059 14679 65117 14680
rect 65163 14720 65205 14729
rect 65163 14680 65164 14720
rect 65204 14680 65205 14720
rect 65163 14671 65205 14680
rect 65355 14720 65397 14729
rect 65355 14680 65356 14720
rect 65396 14680 65397 14720
rect 65355 14671 65397 14680
rect 67939 14720 67997 14721
rect 67939 14680 67948 14720
rect 67988 14680 67997 14720
rect 67939 14679 67997 14680
rect 68803 14720 68861 14721
rect 68803 14680 68812 14720
rect 68852 14680 68861 14720
rect 68803 14679 68861 14680
rect 70347 14720 70389 14729
rect 70347 14680 70348 14720
rect 70388 14680 70389 14720
rect 70347 14671 70389 14680
rect 70723 14720 70781 14721
rect 70723 14680 70732 14720
rect 70772 14680 70781 14720
rect 70723 14679 70781 14680
rect 71587 14720 71645 14721
rect 71587 14680 71596 14720
rect 71636 14680 71645 14720
rect 71587 14679 71645 14680
rect 73611 14720 73653 14729
rect 73611 14680 73612 14720
rect 73652 14680 73653 14720
rect 73611 14671 73653 14680
rect 73803 14720 73845 14729
rect 73803 14680 73804 14720
rect 73844 14680 73845 14720
rect 73803 14671 73845 14680
rect 73891 14720 73949 14721
rect 73891 14680 73900 14720
rect 73940 14680 73949 14720
rect 73891 14679 73949 14680
rect 74091 14720 74133 14729
rect 74091 14680 74092 14720
rect 74132 14680 74133 14720
rect 74091 14671 74133 14680
rect 74187 14720 74229 14729
rect 74187 14680 74188 14720
rect 74228 14680 74229 14720
rect 74187 14671 74229 14680
rect 74283 14720 74325 14729
rect 74283 14680 74284 14720
rect 74324 14680 74325 14720
rect 74283 14671 74325 14680
rect 74379 14720 74421 14729
rect 74379 14680 74380 14720
rect 74420 14680 74421 14720
rect 74379 14671 74421 14680
rect 74659 14720 74717 14721
rect 74659 14680 74668 14720
rect 74708 14680 74717 14720
rect 74659 14679 74717 14680
rect 74955 14720 74997 14729
rect 74955 14680 74956 14720
rect 74996 14680 74997 14720
rect 74955 14671 74997 14680
rect 75627 14720 75669 14729
rect 75627 14680 75628 14720
rect 75668 14680 75669 14720
rect 75627 14671 75669 14680
rect 75819 14720 75861 14729
rect 75819 14680 75820 14720
rect 75860 14680 75861 14720
rect 75819 14671 75861 14680
rect 75907 14720 75965 14721
rect 75907 14680 75916 14720
rect 75956 14680 75965 14720
rect 75907 14679 75965 14680
rect 76203 14720 76245 14729
rect 76203 14680 76204 14720
rect 76244 14680 76245 14720
rect 76203 14671 76245 14680
rect 76579 14720 76637 14721
rect 76579 14680 76588 14720
rect 76628 14680 76637 14720
rect 76579 14679 76637 14680
rect 77443 14720 77501 14721
rect 77443 14680 77452 14720
rect 77492 14680 77501 14720
rect 77443 14679 77501 14680
rect 33003 14650 33045 14659
rect 5163 14636 5205 14645
rect 5163 14596 5164 14636
rect 5204 14596 5205 14636
rect 5163 14587 5205 14596
rect 29931 14636 29973 14645
rect 29931 14596 29932 14636
rect 29972 14596 29973 14636
rect 29931 14587 29973 14596
rect 47499 14636 47541 14645
rect 47499 14596 47500 14636
rect 47540 14596 47541 14636
rect 47499 14587 47541 14596
rect 47979 14636 48021 14645
rect 47979 14596 47980 14636
rect 48020 14596 48021 14636
rect 47979 14587 48021 14596
rect 50763 14636 50805 14645
rect 50763 14596 50764 14636
rect 50804 14596 50805 14636
rect 50763 14587 50805 14596
rect 56427 14636 56469 14645
rect 56427 14596 56428 14636
rect 56468 14596 56469 14636
rect 56427 14587 56469 14596
rect 64395 14636 64437 14645
rect 64395 14596 64396 14636
rect 64436 14596 64437 14636
rect 64395 14587 64437 14596
rect 67563 14636 67605 14645
rect 67563 14596 67564 14636
rect 67604 14596 67605 14636
rect 67563 14587 67605 14596
rect 75051 14636 75093 14645
rect 75051 14596 75052 14636
rect 75092 14596 75093 14636
rect 75051 14587 75093 14596
rect 75723 14636 75765 14645
rect 75723 14596 75724 14636
rect 75764 14596 75765 14636
rect 75723 14587 75765 14596
rect 1035 14552 1077 14561
rect 1035 14512 1036 14552
rect 1076 14512 1077 14552
rect 1035 14503 1077 14512
rect 32323 14552 32381 14553
rect 32323 14512 32332 14552
rect 32372 14512 32381 14552
rect 32323 14511 32381 14512
rect 32707 14552 32765 14553
rect 32707 14512 32716 14552
rect 32756 14512 32765 14552
rect 32707 14511 32765 14512
rect 37411 14552 37469 14553
rect 37411 14512 37420 14552
rect 37460 14512 37469 14552
rect 37411 14511 37469 14512
rect 41539 14552 41597 14553
rect 41539 14512 41548 14552
rect 41588 14512 41597 14552
rect 41539 14511 41597 14512
rect 42883 14552 42941 14553
rect 42883 14512 42892 14552
rect 42932 14512 42941 14552
rect 42883 14511 42941 14512
rect 53155 14552 53213 14553
rect 53155 14512 53164 14552
rect 53204 14512 53213 14552
rect 53155 14511 53213 14512
rect 60555 14552 60597 14561
rect 60555 14512 60556 14552
rect 60596 14512 60597 14552
rect 60555 14503 60597 14512
rect 61803 14552 61845 14561
rect 61803 14512 61804 14552
rect 61844 14512 61845 14552
rect 61803 14503 61845 14512
rect 62571 14552 62613 14561
rect 62571 14512 62572 14552
rect 62612 14512 62613 14552
rect 62571 14503 62613 14512
rect 67371 14552 67413 14561
rect 67371 14512 67372 14552
rect 67412 14512 67413 14552
rect 67371 14503 67413 14512
rect 69955 14552 70013 14553
rect 69955 14512 69964 14552
rect 70004 14512 70013 14552
rect 69955 14511 70013 14512
rect 72739 14552 72797 14553
rect 72739 14512 72748 14552
rect 72788 14512 72797 14552
rect 72739 14511 72797 14512
rect 73699 14552 73757 14553
rect 73699 14512 73708 14552
rect 73748 14512 73757 14552
rect 73699 14511 73757 14512
rect 78595 14552 78653 14553
rect 78595 14512 78604 14552
rect 78644 14512 78653 14552
rect 78595 14511 78653 14512
rect 576 14384 79584 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 76352 14384
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76720 14344 79584 14384
rect 576 14320 79584 14344
rect 1131 14216 1173 14225
rect 1131 14176 1132 14216
rect 1172 14176 1173 14216
rect 1131 14167 1173 14176
rect 2379 14216 2421 14225
rect 2379 14176 2380 14216
rect 2420 14176 2421 14216
rect 2379 14167 2421 14176
rect 2851 14216 2909 14217
rect 2851 14176 2860 14216
rect 2900 14176 2909 14216
rect 2851 14175 2909 14176
rect 7459 14216 7517 14217
rect 7459 14176 7468 14216
rect 7508 14176 7517 14216
rect 7459 14175 7517 14176
rect 35395 14216 35453 14217
rect 35395 14176 35404 14216
rect 35444 14176 35453 14216
rect 35395 14175 35453 14176
rect 38371 14216 38429 14217
rect 38371 14176 38380 14216
rect 38420 14176 38429 14216
rect 38371 14175 38429 14176
rect 39427 14216 39485 14217
rect 39427 14176 39436 14216
rect 39476 14176 39485 14216
rect 39427 14175 39485 14176
rect 51331 14216 51389 14217
rect 51331 14176 51340 14216
rect 51380 14176 51389 14216
rect 51331 14175 51389 14176
rect 52107 14216 52149 14225
rect 52107 14176 52108 14216
rect 52148 14176 52149 14216
rect 52107 14167 52149 14176
rect 56227 14216 56285 14217
rect 56227 14176 56236 14216
rect 56276 14176 56285 14216
rect 56227 14175 56285 14176
rect 68515 14216 68573 14217
rect 68515 14176 68524 14216
rect 68564 14176 68573 14216
rect 68515 14175 68573 14176
rect 69003 14216 69045 14225
rect 69003 14176 69004 14216
rect 69044 14176 69045 14216
rect 69003 14167 69045 14176
rect 70539 14216 70581 14225
rect 70539 14176 70540 14216
rect 70580 14176 70581 14216
rect 70539 14167 70581 14176
rect 79363 14216 79421 14217
rect 79363 14176 79372 14216
rect 79412 14176 79421 14216
rect 79363 14175 79421 14176
rect 32331 14132 32373 14141
rect 32331 14092 32332 14132
rect 32372 14092 32373 14132
rect 32331 14083 32373 14092
rect 40011 14132 40053 14141
rect 40011 14092 40012 14132
rect 40052 14092 40053 14132
rect 40011 14083 40053 14092
rect 43179 14132 43221 14141
rect 43179 14092 43180 14132
rect 43220 14092 43221 14132
rect 43179 14083 43221 14092
rect 47691 14132 47733 14141
rect 47691 14092 47692 14132
rect 47732 14092 47733 14132
rect 47691 14083 47733 14092
rect 52971 14132 53013 14141
rect 52971 14092 52972 14132
rect 53012 14092 53013 14132
rect 52971 14083 53013 14092
rect 68235 14132 68277 14141
rect 68235 14092 68236 14132
rect 68276 14092 68277 14132
rect 70059 14132 70101 14141
rect 68235 14083 68277 14092
rect 68331 14090 68373 14099
rect 2763 14048 2805 14057
rect 2763 14008 2764 14048
rect 2804 14008 2805 14048
rect 2763 13999 2805 14008
rect 2955 14048 2997 14057
rect 2955 14008 2956 14048
rect 2996 14008 2997 14048
rect 2955 13999 2997 14008
rect 3043 14048 3101 14049
rect 3043 14008 3052 14048
rect 3092 14008 3101 14048
rect 3043 14007 3101 14008
rect 4003 14048 4061 14049
rect 4003 14008 4012 14048
rect 4052 14008 4061 14048
rect 4003 14007 4061 14008
rect 4299 14048 4341 14057
rect 4299 14008 4300 14048
rect 4340 14008 4341 14048
rect 4299 13999 4341 14008
rect 4395 14048 4437 14057
rect 4395 14008 4396 14048
rect 4436 14008 4437 14048
rect 4395 13999 4437 14008
rect 5067 14048 5109 14057
rect 5067 14008 5068 14048
rect 5108 14008 5109 14048
rect 5067 13999 5109 14008
rect 5443 14048 5501 14049
rect 5443 14008 5452 14048
rect 5492 14008 5501 14048
rect 5443 14007 5501 14008
rect 6307 14048 6365 14049
rect 6307 14008 6316 14048
rect 6356 14008 6365 14048
rect 6307 14007 6365 14008
rect 31467 14048 31509 14057
rect 31467 14008 31468 14048
rect 31508 14008 31509 14048
rect 31467 13999 31509 14008
rect 31659 14048 31701 14057
rect 31659 14008 31660 14048
rect 31700 14008 31701 14048
rect 31659 13999 31701 14008
rect 31747 14048 31805 14049
rect 31747 14008 31756 14048
rect 31796 14008 31805 14048
rect 31747 14007 31805 14008
rect 32427 14048 32469 14057
rect 32427 14008 32428 14048
rect 32468 14008 32469 14048
rect 32427 13999 32469 14008
rect 32707 14048 32765 14049
rect 32707 14008 32716 14048
rect 32756 14008 32765 14048
rect 32707 14007 32765 14008
rect 33003 14048 33045 14057
rect 33003 14008 33004 14048
rect 33044 14008 33045 14048
rect 33003 13999 33045 14008
rect 33379 14048 33437 14049
rect 33379 14008 33388 14048
rect 33428 14008 33437 14048
rect 33379 14007 33437 14008
rect 34243 14048 34301 14049
rect 34243 14008 34252 14048
rect 34292 14008 34301 14048
rect 34243 14007 34301 14008
rect 37227 14048 37269 14057
rect 37227 14008 37228 14048
rect 37268 14008 37269 14048
rect 37227 13999 37269 14008
rect 38083 14048 38141 14049
rect 38083 14008 38092 14048
rect 38132 14008 38141 14048
rect 38083 14007 38141 14008
rect 38283 14048 38325 14057
rect 38283 14008 38284 14048
rect 38324 14008 38325 14048
rect 38283 13999 38325 14008
rect 38475 14048 38517 14057
rect 38475 14008 38476 14048
rect 38516 14008 38517 14048
rect 38475 13999 38517 14008
rect 38563 14048 38621 14049
rect 38563 14008 38572 14048
rect 38612 14008 38621 14048
rect 38563 14007 38621 14008
rect 39147 14048 39189 14057
rect 39147 14008 39148 14048
rect 39188 14008 39189 14048
rect 39147 13999 39189 14008
rect 39243 14048 39285 14057
rect 39243 14008 39244 14048
rect 39284 14008 39285 14048
rect 39243 13999 39285 14008
rect 39339 14048 39381 14057
rect 39339 14008 39340 14048
rect 39380 14008 39381 14048
rect 39339 13999 39381 14008
rect 39811 14048 39869 14049
rect 39811 14008 39820 14048
rect 39860 14008 39869 14048
rect 39811 14007 39869 14008
rect 39915 14048 39957 14057
rect 39915 14008 39916 14048
rect 39956 14008 39957 14048
rect 39915 13999 39957 14008
rect 40107 14048 40149 14057
rect 40107 14008 40108 14048
rect 40148 14008 40149 14048
rect 40107 13999 40149 14008
rect 40299 14048 40341 14057
rect 40299 14008 40300 14048
rect 40340 14008 40341 14048
rect 40299 13999 40341 14008
rect 40675 14048 40733 14049
rect 40675 14008 40684 14048
rect 40724 14008 40733 14048
rect 40675 14007 40733 14008
rect 41539 14048 41597 14049
rect 41539 14008 41548 14048
rect 41588 14008 41597 14048
rect 41539 14007 41597 14008
rect 43275 14048 43317 14057
rect 43275 14008 43276 14048
rect 43316 14008 43317 14048
rect 43275 13999 43317 14008
rect 43555 14048 43613 14049
rect 43555 14008 43564 14048
rect 43604 14008 43613 14048
rect 43555 14007 43613 14008
rect 44619 14048 44661 14057
rect 44619 14008 44620 14048
rect 44660 14008 44661 14048
rect 44619 13999 44661 14008
rect 44995 14048 45053 14049
rect 44995 14008 45004 14048
rect 45044 14008 45053 14048
rect 44995 14007 45053 14008
rect 45859 14048 45917 14049
rect 45859 14008 45868 14048
rect 45908 14008 45917 14048
rect 45859 14007 45917 14008
rect 47595 14048 47637 14057
rect 47595 14008 47596 14048
rect 47636 14008 47637 14048
rect 47595 13999 47637 14008
rect 47787 14048 47829 14057
rect 47787 14008 47788 14048
rect 47828 14008 47829 14048
rect 47787 13999 47829 14008
rect 47875 14048 47933 14049
rect 47875 14008 47884 14048
rect 47924 14008 47933 14048
rect 47875 14007 47933 14008
rect 51139 14048 51197 14049
rect 51139 14008 51148 14048
rect 51188 14008 51197 14048
rect 51139 14007 51197 14008
rect 51243 14048 51285 14057
rect 51243 14008 51244 14048
rect 51284 14008 51285 14048
rect 51243 13999 51285 14008
rect 51435 14048 51477 14057
rect 51435 14008 51436 14048
rect 51476 14008 51477 14048
rect 51435 13999 51477 14008
rect 52579 14048 52637 14049
rect 52579 14008 52588 14048
rect 52628 14008 52637 14048
rect 52579 14007 52637 14008
rect 52875 14048 52917 14057
rect 52875 14008 52876 14048
rect 52916 14008 52917 14048
rect 52875 13999 52917 14008
rect 53059 14048 53117 14049
rect 53059 14008 53068 14048
rect 53108 14008 53117 14048
rect 53059 14007 53117 14008
rect 53347 14048 53405 14049
rect 53347 14008 53356 14048
rect 53396 14008 53405 14048
rect 53347 14007 53405 14008
rect 53451 14048 53493 14057
rect 53451 14008 53452 14048
rect 53492 14008 53493 14048
rect 53451 13999 53493 14008
rect 53643 14048 53685 14057
rect 53643 14008 53644 14048
rect 53684 14008 53685 14048
rect 53643 13999 53685 14008
rect 53835 14048 53877 14057
rect 53835 14008 53836 14048
rect 53876 14008 53877 14048
rect 53835 13999 53877 14008
rect 54211 14048 54269 14049
rect 54211 14008 54220 14048
rect 54260 14008 54269 14048
rect 54211 14007 54269 14008
rect 55075 14048 55133 14049
rect 55075 14008 55084 14048
rect 55124 14008 55133 14048
rect 55075 14007 55133 14008
rect 56419 14048 56477 14049
rect 56419 14008 56428 14048
rect 56468 14008 56477 14048
rect 56419 14007 56477 14008
rect 56619 14048 56661 14057
rect 56619 14008 56620 14048
rect 56660 14008 56661 14048
rect 56619 13999 56661 14008
rect 57763 14048 57821 14049
rect 57763 14008 57772 14048
rect 57812 14008 57821 14048
rect 57763 14007 57821 14008
rect 57963 14048 58005 14057
rect 57963 14008 57964 14048
rect 58004 14008 58005 14048
rect 57963 13999 58005 14008
rect 58155 14048 58197 14057
rect 58155 14008 58156 14048
rect 58196 14008 58197 14048
rect 58155 13999 58197 14008
rect 58531 14048 58589 14049
rect 58531 14008 58540 14048
rect 58580 14008 58589 14048
rect 58531 14007 58589 14008
rect 59395 14048 59453 14049
rect 59395 14008 59404 14048
rect 59444 14008 59453 14048
rect 59395 14007 59453 14008
rect 60835 14048 60893 14049
rect 60835 14008 60844 14048
rect 60884 14008 60893 14048
rect 60835 14007 60893 14008
rect 61035 14048 61077 14057
rect 61035 14008 61036 14048
rect 61076 14008 61077 14048
rect 61035 13999 61077 14008
rect 61227 14048 61269 14057
rect 61227 14008 61228 14048
rect 61268 14008 61269 14048
rect 61227 13999 61269 14008
rect 61603 14048 61661 14049
rect 61603 14008 61612 14048
rect 61652 14008 61661 14048
rect 61603 14007 61661 14008
rect 62467 14048 62525 14049
rect 62467 14008 62476 14048
rect 62516 14008 62525 14048
rect 62467 14007 62525 14008
rect 63811 14048 63869 14049
rect 63811 14008 63820 14048
rect 63860 14008 63869 14048
rect 63811 14007 63869 14008
rect 63915 14048 63957 14057
rect 63915 14008 63916 14048
rect 63956 14008 63957 14048
rect 63915 13999 63957 14008
rect 64107 14048 64149 14057
rect 64107 14008 64108 14048
rect 64148 14008 64149 14048
rect 64107 13999 64149 14008
rect 64683 14048 64725 14057
rect 64683 14008 64684 14048
rect 64724 14008 64725 14048
rect 64683 13999 64725 14008
rect 65059 14048 65117 14049
rect 65059 14008 65068 14048
rect 65108 14008 65117 14048
rect 65059 14007 65117 14008
rect 65923 14048 65981 14049
rect 65923 14008 65932 14048
rect 65972 14008 65981 14048
rect 65923 14007 65981 14008
rect 67267 14048 67325 14049
rect 67267 14008 67276 14048
rect 67316 14008 67325 14048
rect 67267 14007 67325 14008
rect 67371 14048 67413 14057
rect 67371 14008 67372 14048
rect 67412 14008 67413 14048
rect 67371 13999 67413 14008
rect 67563 14048 67605 14057
rect 67563 14008 67564 14048
rect 67604 14008 67605 14048
rect 67563 13999 67605 14008
rect 68035 14048 68093 14049
rect 68035 14008 68044 14048
rect 68084 14008 68093 14048
rect 68035 14007 68093 14008
rect 68139 14048 68181 14057
rect 68139 14008 68140 14048
rect 68180 14008 68181 14048
rect 68331 14050 68332 14090
rect 68372 14050 68373 14090
rect 70059 14092 70060 14132
rect 70100 14092 70101 14132
rect 70059 14083 70101 14092
rect 71019 14132 71061 14141
rect 71019 14092 71020 14132
rect 71060 14092 71061 14132
rect 71019 14083 71061 14092
rect 72171 14132 72213 14141
rect 72171 14092 72172 14132
rect 72212 14092 72213 14132
rect 72171 14083 72213 14092
rect 75915 14132 75957 14141
rect 75915 14092 75916 14132
rect 75956 14092 75957 14132
rect 75915 14083 75957 14092
rect 68331 14041 68373 14050
rect 68619 14069 68661 14078
rect 68619 14029 68620 14069
rect 68660 14029 68661 14069
rect 68619 14020 68661 14029
rect 68715 14048 68757 14057
rect 68139 13999 68181 14008
rect 68715 14008 68716 14048
rect 68756 14008 68757 14048
rect 68715 13999 68757 14008
rect 68811 14048 68853 14057
rect 68811 14008 68812 14048
rect 68852 14008 68853 14048
rect 68811 13999 68853 14008
rect 69667 14048 69725 14049
rect 69667 14008 69676 14048
rect 69716 14008 69725 14048
rect 69667 14007 69725 14008
rect 69963 14048 70005 14057
rect 69963 14008 69964 14048
rect 70004 14008 70005 14048
rect 69963 13999 70005 14008
rect 70915 14048 70973 14049
rect 70915 14008 70924 14048
rect 70964 14008 70973 14048
rect 70915 14007 70973 14008
rect 71115 14048 71157 14057
rect 71115 14008 71116 14048
rect 71156 14008 71157 14048
rect 71115 13999 71157 14008
rect 72547 14048 72605 14049
rect 72547 14008 72556 14048
rect 72596 14008 72605 14048
rect 74763 14048 74805 14057
rect 72547 14007 72605 14008
rect 73411 14037 73469 14038
rect 73411 13997 73420 14037
rect 73460 13997 73469 14037
rect 74763 14008 74764 14048
rect 74804 14008 74805 14048
rect 74763 13999 74805 14008
rect 74955 14048 74997 14057
rect 74955 14008 74956 14048
rect 74996 14008 74997 14048
rect 74955 13999 74997 14008
rect 75043 14048 75101 14049
rect 75043 14008 75052 14048
rect 75092 14008 75101 14048
rect 75043 14007 75101 14008
rect 75811 14048 75869 14049
rect 75811 14008 75820 14048
rect 75860 14008 75869 14048
rect 75811 14007 75869 14008
rect 76011 14048 76053 14057
rect 76011 14008 76012 14048
rect 76052 14008 76053 14048
rect 76011 13999 76053 14008
rect 76971 14048 77013 14057
rect 76971 14008 76972 14048
rect 77012 14008 77013 14048
rect 76971 13999 77013 14008
rect 77347 14048 77405 14049
rect 77347 14008 77356 14048
rect 77396 14008 77405 14048
rect 77347 14007 77405 14008
rect 78211 14048 78269 14049
rect 78211 14008 78220 14048
rect 78260 14008 78269 14048
rect 78211 14007 78269 14008
rect 73411 13996 73469 13997
rect 1315 13964 1373 13965
rect 1315 13924 1324 13964
rect 1364 13924 1373 13964
rect 1315 13923 1373 13924
rect 1699 13964 1757 13965
rect 1699 13924 1708 13964
rect 1748 13924 1757 13964
rect 1699 13923 1757 13924
rect 2563 13964 2621 13965
rect 2563 13924 2572 13964
rect 2612 13924 2621 13964
rect 2563 13923 2621 13924
rect 47019 13964 47061 13973
rect 47019 13924 47020 13964
rect 47060 13924 47061 13964
rect 47019 13915 47061 13924
rect 67083 13964 67125 13973
rect 67083 13924 67084 13964
rect 67124 13924 67125 13964
rect 67083 13915 67125 13924
rect 69187 13964 69245 13965
rect 69187 13924 69196 13964
rect 69236 13924 69245 13964
rect 69187 13923 69245 13924
rect 70723 13964 70781 13965
rect 70723 13924 70732 13964
rect 70772 13924 70781 13964
rect 70723 13923 70781 13924
rect 30411 13880 30453 13889
rect 30411 13840 30412 13880
rect 30452 13840 30453 13880
rect 30411 13831 30453 13840
rect 31467 13880 31509 13889
rect 31467 13840 31468 13880
rect 31508 13840 31509 13880
rect 31467 13831 31509 13840
rect 43851 13880 43893 13889
rect 43851 13840 43852 13880
rect 43892 13840 43893 13880
rect 43851 13831 43893 13840
rect 50955 13880 50997 13889
rect 50955 13840 50956 13880
rect 50996 13840 50997 13880
rect 50955 13831 50997 13840
rect 67563 13880 67605 13889
rect 67563 13840 67564 13880
rect 67604 13840 67605 13880
rect 67563 13831 67605 13840
rect 1515 13796 1557 13805
rect 1515 13756 1516 13796
rect 1556 13756 1557 13796
rect 1515 13747 1557 13756
rect 4675 13796 4733 13797
rect 4675 13756 4684 13796
rect 4724 13756 4733 13796
rect 4675 13755 4733 13756
rect 32035 13796 32093 13797
rect 32035 13756 32044 13796
rect 32084 13756 32093 13796
rect 32035 13755 32093 13756
rect 37611 13796 37653 13805
rect 37611 13756 37612 13796
rect 37652 13756 37653 13796
rect 37611 13747 37653 13756
rect 42691 13796 42749 13797
rect 42691 13756 42700 13796
rect 42740 13756 42749 13796
rect 42691 13755 42749 13756
rect 42883 13796 42941 13797
rect 42883 13756 42892 13796
rect 42932 13756 42941 13796
rect 42883 13755 42941 13756
rect 53643 13796 53685 13805
rect 53643 13756 53644 13796
rect 53684 13756 53685 13796
rect 53643 13747 53685 13756
rect 56227 13796 56285 13797
rect 56227 13756 56236 13796
rect 56276 13756 56285 13796
rect 56227 13755 56285 13756
rect 56523 13796 56565 13805
rect 56523 13756 56524 13796
rect 56564 13756 56565 13796
rect 56523 13747 56565 13756
rect 57867 13796 57909 13805
rect 57867 13756 57868 13796
rect 57908 13756 57909 13796
rect 57867 13747 57909 13756
rect 60547 13796 60605 13797
rect 60547 13756 60556 13796
rect 60596 13756 60605 13796
rect 60547 13755 60605 13756
rect 60939 13796 60981 13805
rect 60939 13756 60940 13796
rect 60980 13756 60981 13796
rect 60939 13747 60981 13756
rect 63619 13796 63677 13797
rect 63619 13756 63628 13796
rect 63668 13756 63677 13796
rect 63619 13755 63677 13756
rect 64107 13796 64149 13805
rect 64107 13756 64108 13796
rect 64148 13756 64149 13796
rect 64107 13747 64149 13756
rect 70339 13796 70397 13797
rect 70339 13756 70348 13796
rect 70388 13756 70397 13796
rect 70339 13755 70397 13756
rect 74563 13796 74621 13797
rect 74563 13756 74572 13796
rect 74612 13756 74621 13796
rect 74563 13755 74621 13756
rect 74763 13796 74805 13805
rect 74763 13756 74764 13796
rect 74804 13756 74805 13796
rect 74763 13747 74805 13756
rect 576 13628 79584 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 75112 13628
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75480 13588 79584 13628
rect 576 13564 79584 13588
rect 4483 13460 4541 13461
rect 4483 13420 4492 13460
rect 4532 13420 4541 13460
rect 4483 13419 4541 13420
rect 32427 13460 32469 13469
rect 32427 13420 32428 13460
rect 32468 13420 32469 13460
rect 32427 13411 32469 13420
rect 33003 13460 33045 13469
rect 33003 13420 33004 13460
rect 33044 13420 33045 13460
rect 33003 13411 33045 13420
rect 36267 13460 36309 13469
rect 36267 13420 36268 13460
rect 36308 13420 36309 13460
rect 36267 13411 36309 13420
rect 41547 13460 41589 13469
rect 41547 13420 41548 13460
rect 41588 13420 41589 13460
rect 41547 13411 41589 13420
rect 42795 13460 42837 13469
rect 42795 13420 42796 13460
rect 42836 13420 42837 13460
rect 42795 13411 42837 13420
rect 45475 13460 45533 13461
rect 45475 13420 45484 13460
rect 45524 13420 45533 13460
rect 45475 13419 45533 13420
rect 47307 13460 47349 13469
rect 47307 13420 47308 13460
rect 47348 13420 47349 13460
rect 47307 13411 47349 13420
rect 54699 13460 54741 13469
rect 54699 13420 54700 13460
rect 54740 13420 54741 13460
rect 54699 13411 54741 13420
rect 58731 13460 58773 13469
rect 58731 13420 58732 13460
rect 58772 13420 58773 13460
rect 58731 13411 58773 13420
rect 61027 13460 61085 13461
rect 61027 13420 61036 13460
rect 61076 13420 61085 13460
rect 61027 13419 61085 13420
rect 64587 13460 64629 13469
rect 64587 13420 64588 13460
rect 64628 13420 64629 13460
rect 64587 13411 64629 13420
rect 70155 13460 70197 13469
rect 70155 13420 70156 13460
rect 70196 13420 70197 13460
rect 70155 13411 70197 13420
rect 76491 13460 76533 13469
rect 76491 13420 76492 13460
rect 76532 13420 76533 13460
rect 76491 13411 76533 13420
rect 1227 13376 1269 13385
rect 1227 13336 1228 13376
rect 1268 13336 1269 13376
rect 1227 13327 1269 13336
rect 1899 13376 1941 13385
rect 1899 13336 1900 13376
rect 1940 13336 1941 13376
rect 1899 13327 1941 13336
rect 5355 13376 5397 13385
rect 5355 13336 5356 13376
rect 5396 13336 5397 13376
rect 5355 13327 5397 13336
rect 6219 13376 6261 13385
rect 6219 13336 6220 13376
rect 6260 13336 6261 13376
rect 6219 13327 6261 13336
rect 39531 13376 39573 13385
rect 39531 13336 39532 13376
rect 39572 13336 39573 13376
rect 39531 13327 39573 13336
rect 40779 13376 40821 13385
rect 40779 13336 40780 13376
rect 40820 13336 40821 13376
rect 40779 13327 40821 13336
rect 51811 13376 51869 13377
rect 51811 13336 51820 13376
rect 51860 13336 51869 13376
rect 51811 13335 51869 13336
rect 56331 13376 56373 13385
rect 56331 13336 56332 13376
rect 56372 13336 56373 13376
rect 56331 13327 56373 13336
rect 58531 13376 58589 13377
rect 58531 13336 58540 13376
rect 58580 13336 58589 13376
rect 58531 13335 58589 13336
rect 62475 13376 62517 13385
rect 62475 13336 62476 13376
rect 62516 13336 62517 13376
rect 62475 13327 62517 13336
rect 65163 13376 65205 13385
rect 65163 13336 65164 13376
rect 65204 13336 65205 13376
rect 65163 13327 65205 13336
rect 71019 13376 71061 13385
rect 71019 13336 71020 13376
rect 71060 13336 71061 13376
rect 71019 13327 71061 13336
rect 71979 13376 72021 13385
rect 71979 13336 71980 13376
rect 72020 13336 72021 13376
rect 71979 13327 72021 13336
rect 74563 13376 74621 13377
rect 74563 13336 74572 13376
rect 74612 13336 74621 13376
rect 74563 13335 74621 13336
rect 76099 13376 76157 13377
rect 76099 13336 76108 13376
rect 76148 13336 76157 13376
rect 76099 13335 76157 13336
rect 77067 13376 77109 13385
rect 77067 13336 77068 13376
rect 77108 13336 77109 13376
rect 77067 13327 77109 13336
rect 77451 13376 77493 13385
rect 77451 13336 77452 13376
rect 77492 13336 77493 13376
rect 77451 13327 77493 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1411 13292 1469 13293
rect 1411 13252 1420 13292
rect 1460 13252 1469 13292
rect 1411 13251 1469 13252
rect 6699 13292 6741 13301
rect 6699 13252 6700 13292
rect 6740 13252 6741 13292
rect 6699 13243 6741 13252
rect 48067 13250 48125 13251
rect 36163 13231 36221 13232
rect 1603 13208 1661 13209
rect 1603 13168 1612 13208
rect 1652 13168 1661 13208
rect 1603 13167 1661 13168
rect 1707 13208 1749 13217
rect 1707 13168 1708 13208
rect 1748 13168 1749 13208
rect 1707 13159 1749 13168
rect 1899 13208 1941 13217
rect 1899 13168 1900 13208
rect 1940 13168 1941 13208
rect 1899 13159 1941 13168
rect 2091 13208 2133 13217
rect 2091 13168 2092 13208
rect 2132 13168 2133 13208
rect 2091 13159 2133 13168
rect 2467 13208 2525 13209
rect 2467 13168 2476 13208
rect 2516 13168 2525 13208
rect 2467 13167 2525 13168
rect 3331 13208 3389 13209
rect 3331 13168 3340 13208
rect 3380 13168 3389 13208
rect 3331 13167 3389 13168
rect 5163 13208 5205 13217
rect 5163 13168 5164 13208
rect 5204 13168 5205 13208
rect 5163 13159 5205 13168
rect 6019 13208 6077 13209
rect 6019 13168 6028 13208
rect 6068 13168 6077 13208
rect 6019 13167 6077 13168
rect 6603 13208 6645 13217
rect 6603 13168 6604 13208
rect 6644 13168 6645 13208
rect 6603 13159 6645 13168
rect 6787 13208 6845 13209
rect 6787 13168 6796 13208
rect 6836 13168 6845 13208
rect 6787 13167 6845 13168
rect 32331 13208 32373 13217
rect 32331 13168 32332 13208
rect 32372 13168 32373 13208
rect 32331 13159 32373 13168
rect 32515 13208 32573 13209
rect 32515 13168 32524 13208
rect 32564 13168 32573 13208
rect 32515 13167 32573 13168
rect 32707 13208 32765 13209
rect 32707 13168 32716 13208
rect 32756 13168 32765 13208
rect 32707 13167 32765 13168
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 33003 13208 33045 13217
rect 33003 13168 33004 13208
rect 33044 13168 33045 13208
rect 33003 13159 33045 13168
rect 34819 13208 34877 13209
rect 34819 13168 34828 13208
rect 34868 13168 34877 13208
rect 34819 13167 34877 13168
rect 34923 13208 34965 13217
rect 34923 13168 34924 13208
rect 34964 13168 34965 13208
rect 34923 13159 34965 13168
rect 35115 13208 35157 13217
rect 35115 13168 35116 13208
rect 35156 13168 35157 13208
rect 36163 13191 36172 13231
rect 36212 13191 36221 13231
rect 47491 13222 47549 13223
rect 36163 13190 36221 13191
rect 36363 13208 36405 13217
rect 35115 13159 35157 13168
rect 36363 13168 36364 13208
rect 36404 13168 36405 13208
rect 36363 13159 36405 13168
rect 36547 13208 36605 13209
rect 36547 13168 36556 13208
rect 36596 13168 36605 13208
rect 36547 13167 36605 13168
rect 36747 13208 36789 13217
rect 36747 13168 36748 13208
rect 36788 13168 36789 13208
rect 36747 13159 36789 13168
rect 37315 13208 37373 13209
rect 37315 13168 37324 13208
rect 37364 13168 37373 13208
rect 37315 13167 37373 13168
rect 38179 13208 38237 13209
rect 38179 13168 38188 13208
rect 38228 13168 38237 13208
rect 38179 13167 38237 13168
rect 41547 13208 41589 13217
rect 41547 13168 41548 13208
rect 41588 13168 41589 13208
rect 41547 13159 41589 13168
rect 41739 13208 41781 13217
rect 41739 13168 41740 13208
rect 41780 13168 41781 13208
rect 41739 13159 41781 13168
rect 41827 13208 41885 13209
rect 41827 13168 41836 13208
rect 41876 13168 41885 13208
rect 41827 13167 41885 13168
rect 42691 13208 42749 13209
rect 42691 13168 42700 13208
rect 42740 13168 42749 13208
rect 42691 13167 42749 13168
rect 42891 13208 42933 13217
rect 42891 13168 42892 13208
rect 42932 13168 42933 13208
rect 42891 13159 42933 13168
rect 43083 13208 43125 13217
rect 43083 13168 43084 13208
rect 43124 13168 43125 13208
rect 43083 13159 43125 13168
rect 43459 13208 43517 13209
rect 43459 13168 43468 13208
rect 43508 13168 43517 13208
rect 43459 13167 43517 13168
rect 44323 13208 44381 13209
rect 44323 13168 44332 13208
rect 44372 13168 44381 13208
rect 44323 13167 44381 13168
rect 46147 13208 46205 13209
rect 46147 13168 46156 13208
rect 46196 13168 46205 13208
rect 46147 13167 46205 13168
rect 47307 13208 47349 13217
rect 47307 13168 47308 13208
rect 47348 13168 47349 13208
rect 47491 13182 47500 13222
rect 47540 13182 47549 13222
rect 47491 13181 47549 13182
rect 47587 13208 47645 13209
rect 47307 13159 47349 13168
rect 47587 13168 47596 13208
rect 47636 13168 47645 13208
rect 47587 13167 47645 13168
rect 47883 13208 47925 13217
rect 47883 13168 47884 13208
rect 47924 13168 47925 13208
rect 47883 13159 47925 13168
rect 47979 13208 48021 13217
rect 48067 13210 48076 13250
rect 48116 13210 48125 13250
rect 73411 13219 73469 13220
rect 48067 13209 48125 13210
rect 47979 13168 47980 13208
rect 48020 13168 48021 13208
rect 47979 13159 48021 13168
rect 48643 13208 48701 13209
rect 48643 13168 48652 13208
rect 48692 13168 48701 13208
rect 48643 13167 48701 13168
rect 48843 13208 48885 13217
rect 48843 13168 48844 13208
rect 48884 13168 48885 13208
rect 48843 13159 48885 13168
rect 49795 13208 49853 13209
rect 49795 13168 49804 13208
rect 49844 13168 49853 13208
rect 49795 13167 49853 13168
rect 50659 13208 50717 13209
rect 50659 13168 50668 13208
rect 50708 13168 50717 13208
rect 50659 13167 50717 13168
rect 54403 13208 54461 13209
rect 54403 13168 54412 13208
rect 54452 13168 54461 13208
rect 54403 13167 54461 13168
rect 54507 13208 54549 13217
rect 54507 13168 54508 13208
rect 54548 13168 54549 13208
rect 54507 13159 54549 13168
rect 54699 13208 54741 13217
rect 54699 13168 54700 13208
rect 54740 13168 54741 13208
rect 54699 13159 54741 13168
rect 55083 13208 55125 13217
rect 55083 13168 55084 13208
rect 55124 13168 55125 13208
rect 55083 13159 55125 13168
rect 55179 13208 55221 13217
rect 55179 13168 55180 13208
rect 55220 13168 55221 13208
rect 55179 13159 55221 13168
rect 55275 13208 55317 13217
rect 55275 13168 55276 13208
rect 55316 13168 55317 13208
rect 55275 13159 55317 13168
rect 55371 13208 55413 13217
rect 55371 13168 55372 13208
rect 55412 13168 55413 13208
rect 55371 13159 55413 13168
rect 56035 13208 56093 13209
rect 56035 13168 56044 13208
rect 56084 13168 56093 13208
rect 56035 13167 56093 13168
rect 56139 13208 56181 13217
rect 56139 13168 56140 13208
rect 56180 13168 56181 13208
rect 56139 13159 56181 13168
rect 56331 13208 56373 13217
rect 56331 13168 56332 13208
rect 56372 13168 56373 13208
rect 56331 13159 56373 13168
rect 56523 13208 56565 13217
rect 56523 13168 56524 13208
rect 56564 13168 56565 13208
rect 56523 13159 56565 13168
rect 56715 13208 56757 13217
rect 56715 13168 56716 13208
rect 56756 13168 56757 13208
rect 56715 13159 56757 13168
rect 56803 13208 56861 13209
rect 56803 13168 56812 13208
rect 56852 13168 56861 13208
rect 56803 13167 56861 13168
rect 57859 13208 57917 13209
rect 57859 13168 57868 13208
rect 57908 13168 57917 13208
rect 57859 13167 57917 13168
rect 58155 13208 58197 13217
rect 58155 13168 58156 13208
rect 58196 13168 58197 13208
rect 58155 13159 58197 13168
rect 58731 13208 58773 13217
rect 58731 13168 58732 13208
rect 58772 13168 58773 13208
rect 58731 13159 58773 13168
rect 58923 13208 58965 13217
rect 58923 13168 58924 13208
rect 58964 13168 58965 13208
rect 58923 13159 58965 13168
rect 59011 13208 59069 13209
rect 59011 13168 59020 13208
rect 59060 13168 59069 13208
rect 59011 13167 59069 13168
rect 61323 13208 61365 13217
rect 61323 13168 61324 13208
rect 61364 13168 61365 13208
rect 61323 13159 61365 13168
rect 61419 13208 61461 13217
rect 61419 13168 61420 13208
rect 61460 13168 61461 13208
rect 61419 13159 61461 13168
rect 61699 13208 61757 13209
rect 61699 13168 61708 13208
rect 61748 13168 61757 13208
rect 61699 13167 61757 13168
rect 62091 13208 62133 13217
rect 62091 13168 62092 13208
rect 62132 13168 62133 13208
rect 62091 13159 62133 13168
rect 62187 13208 62229 13217
rect 62187 13168 62188 13208
rect 62228 13168 62229 13208
rect 62187 13159 62229 13168
rect 62283 13208 62325 13217
rect 62283 13168 62284 13208
rect 62324 13168 62325 13208
rect 62283 13159 62325 13168
rect 63915 13208 63957 13217
rect 63915 13168 63916 13208
rect 63956 13168 63957 13208
rect 63915 13159 63957 13168
rect 64011 13208 64053 13217
rect 64011 13168 64012 13208
rect 64052 13168 64053 13208
rect 64011 13159 64053 13168
rect 64107 13208 64149 13217
rect 64107 13168 64108 13208
rect 64148 13168 64149 13208
rect 64107 13159 64149 13168
rect 64291 13208 64349 13209
rect 64291 13168 64300 13208
rect 64340 13168 64349 13208
rect 64291 13167 64349 13168
rect 64395 13208 64437 13217
rect 64395 13168 64396 13208
rect 64436 13168 64437 13208
rect 64395 13159 64437 13168
rect 64587 13208 64629 13217
rect 64587 13168 64588 13208
rect 64628 13168 64629 13208
rect 64587 13159 64629 13168
rect 68715 13208 68757 13217
rect 68715 13168 68716 13208
rect 68756 13168 68757 13208
rect 68715 13159 68757 13168
rect 68811 13208 68853 13217
rect 68811 13168 68812 13208
rect 68852 13168 68853 13208
rect 68811 13159 68853 13168
rect 68907 13208 68949 13217
rect 68907 13168 68908 13208
rect 68948 13168 68949 13208
rect 68907 13159 68949 13168
rect 69099 13208 69141 13217
rect 69099 13168 69100 13208
rect 69140 13168 69141 13208
rect 69099 13159 69141 13168
rect 69291 13208 69333 13217
rect 69291 13168 69292 13208
rect 69332 13168 69333 13208
rect 69291 13159 69333 13168
rect 69379 13208 69437 13209
rect 69379 13168 69388 13208
rect 69428 13168 69437 13208
rect 69379 13167 69437 13168
rect 69667 13208 69725 13209
rect 69667 13168 69676 13208
rect 69716 13168 69725 13208
rect 69667 13167 69725 13168
rect 69867 13208 69909 13217
rect 69867 13168 69868 13208
rect 69908 13168 69909 13208
rect 69867 13159 69909 13168
rect 70051 13208 70109 13209
rect 70051 13168 70060 13208
rect 70100 13168 70109 13208
rect 70051 13167 70109 13168
rect 70251 13208 70293 13217
rect 70251 13168 70252 13208
rect 70292 13168 70293 13208
rect 70251 13159 70293 13168
rect 72171 13208 72213 13217
rect 72171 13168 72172 13208
rect 72212 13168 72213 13208
rect 72171 13159 72213 13168
rect 72547 13208 72605 13209
rect 72547 13168 72556 13208
rect 72596 13168 72605 13208
rect 73411 13179 73420 13219
rect 73460 13179 73469 13219
rect 73411 13178 73469 13179
rect 74763 13208 74805 13217
rect 72547 13167 72605 13168
rect 74763 13168 74764 13208
rect 74804 13168 74805 13208
rect 74763 13159 74805 13168
rect 74859 13208 74901 13217
rect 74859 13168 74860 13208
rect 74900 13168 74901 13208
rect 74859 13159 74901 13168
rect 74955 13208 74997 13217
rect 74955 13168 74956 13208
rect 74996 13168 74997 13208
rect 74955 13159 74997 13168
rect 75051 13208 75093 13217
rect 75051 13168 75052 13208
rect 75092 13168 75093 13208
rect 75051 13159 75093 13168
rect 75427 13208 75485 13209
rect 75427 13168 75436 13208
rect 75476 13168 75485 13208
rect 75427 13167 75485 13168
rect 75723 13208 75765 13217
rect 75723 13168 75724 13208
rect 75764 13168 75765 13208
rect 75723 13159 75765 13168
rect 75819 13208 75861 13217
rect 75819 13168 75820 13208
rect 75860 13168 75861 13208
rect 75819 13159 75861 13168
rect 76491 13208 76533 13217
rect 76491 13168 76492 13208
rect 76532 13168 76533 13208
rect 76491 13159 76533 13168
rect 76683 13208 76725 13217
rect 76683 13168 76684 13208
rect 76724 13168 76725 13208
rect 76683 13159 76725 13168
rect 76771 13208 76829 13209
rect 76771 13168 76780 13208
rect 76820 13168 76829 13208
rect 76771 13167 76829 13168
rect 76963 13208 77021 13209
rect 76963 13168 76972 13208
rect 77012 13168 77021 13208
rect 76963 13167 77021 13168
rect 77163 13208 77205 13217
rect 77163 13168 77164 13208
rect 77204 13168 77205 13208
rect 77163 13159 77205 13168
rect 36651 13124 36693 13133
rect 36651 13084 36652 13124
rect 36692 13084 36693 13124
rect 36651 13075 36693 13084
rect 36939 13124 36981 13133
rect 36939 13084 36940 13124
rect 36980 13084 36981 13124
rect 36939 13075 36981 13084
rect 48747 13124 48789 13133
rect 48747 13084 48748 13124
rect 48788 13084 48789 13124
rect 48747 13075 48789 13084
rect 49419 13124 49461 13133
rect 49419 13084 49420 13124
rect 49460 13084 49461 13124
rect 49419 13075 49461 13084
rect 58251 13124 58293 13133
rect 58251 13084 58252 13124
rect 58292 13084 58293 13124
rect 58251 13075 58293 13084
rect 69771 13124 69813 13133
rect 69771 13084 69772 13124
rect 69812 13084 69813 13124
rect 69771 13075 69813 13084
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 35011 13040 35069 13041
rect 35011 13000 35020 13040
rect 35060 13000 35069 13040
rect 35011 12999 35069 13000
rect 39331 13040 39389 13041
rect 39331 13000 39340 13040
rect 39380 13000 39389 13040
rect 39331 12999 39389 13000
rect 46635 13040 46677 13049
rect 46635 13000 46636 13040
rect 46676 13000 46677 13040
rect 46635 12991 46677 13000
rect 48163 13040 48221 13041
rect 48163 13000 48172 13040
rect 48212 13000 48221 13040
rect 48163 12999 48221 13000
rect 56611 13040 56669 13041
rect 56611 13000 56620 13040
rect 56660 13000 56669 13040
rect 56611 12999 56669 13000
rect 61987 13040 62045 13041
rect 61987 13000 61996 13040
rect 62036 13000 62045 13040
rect 61987 12999 62045 13000
rect 63811 13040 63869 13041
rect 63811 13000 63820 13040
rect 63860 13000 63869 13040
rect 63811 12999 63869 13000
rect 68611 13040 68669 13041
rect 68611 13000 68620 13040
rect 68660 13000 68669 13040
rect 68611 12999 68669 13000
rect 69187 13040 69245 13041
rect 69187 13000 69196 13040
rect 69236 13000 69245 13040
rect 69187 12999 69245 13000
rect 576 12872 79584 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 76352 12872
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76720 12832 79584 12872
rect 576 12808 79584 12832
rect 1891 12704 1949 12705
rect 1891 12664 1900 12704
rect 1940 12664 1949 12704
rect 1891 12663 1949 12664
rect 4579 12704 4637 12705
rect 4579 12664 4588 12704
rect 4628 12664 4637 12704
rect 4579 12663 4637 12664
rect 41443 12704 41501 12705
rect 41443 12664 41452 12704
rect 41492 12664 41501 12704
rect 41443 12663 41501 12664
rect 47875 12704 47933 12705
rect 47875 12664 47884 12704
rect 47924 12664 47933 12704
rect 47875 12663 47933 12664
rect 49123 12704 49181 12705
rect 49123 12664 49132 12704
rect 49172 12664 49181 12704
rect 49123 12663 49181 12664
rect 57283 12704 57341 12705
rect 57283 12664 57292 12704
rect 57332 12664 57341 12704
rect 57283 12663 57341 12664
rect 61411 12704 61469 12705
rect 61411 12664 61420 12704
rect 61460 12664 61469 12704
rect 61411 12663 61469 12664
rect 67171 12704 67229 12705
rect 67171 12664 67180 12704
rect 67220 12664 67229 12704
rect 67171 12663 67229 12664
rect 72835 12704 72893 12705
rect 72835 12664 72844 12704
rect 72884 12664 72893 12704
rect 72835 12663 72893 12664
rect 74371 12704 74429 12705
rect 74371 12664 74380 12704
rect 74420 12664 74429 12704
rect 74371 12663 74429 12664
rect 48555 12620 48597 12629
rect 48555 12580 48556 12620
rect 48596 12580 48597 12620
rect 48555 12571 48597 12580
rect 54891 12620 54933 12629
rect 54891 12580 54892 12620
rect 54932 12580 54933 12620
rect 76107 12620 76149 12629
rect 54891 12571 54933 12580
rect 74763 12578 74805 12587
rect 1995 12557 2037 12566
rect 1995 12517 1996 12557
rect 2036 12517 2037 12557
rect 1995 12508 2037 12517
rect 2091 12557 2133 12566
rect 2091 12517 2092 12557
rect 2132 12517 2133 12557
rect 2091 12508 2133 12517
rect 2379 12536 2421 12545
rect 2187 12491 2229 12500
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1315 12452 1373 12453
rect 1315 12412 1324 12452
rect 1364 12412 1373 12452
rect 1315 12411 1373 12412
rect 1699 12452 1757 12453
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 2187 12451 2188 12491
rect 2228 12451 2229 12491
rect 2379 12496 2380 12536
rect 2420 12496 2421 12536
rect 2379 12487 2421 12496
rect 2571 12536 2613 12545
rect 2571 12496 2572 12536
rect 2612 12496 2613 12536
rect 2571 12487 2613 12496
rect 2659 12536 2717 12537
rect 2659 12496 2668 12536
rect 2708 12496 2717 12536
rect 2659 12495 2717 12496
rect 4491 12536 4533 12545
rect 4491 12496 4492 12536
rect 4532 12496 4533 12536
rect 4491 12487 4533 12496
rect 4683 12536 4725 12545
rect 4683 12496 4684 12536
rect 4724 12496 4725 12536
rect 4683 12487 4725 12496
rect 4771 12536 4829 12537
rect 4771 12496 4780 12536
rect 4820 12496 4829 12536
rect 4771 12495 4829 12496
rect 5355 12536 5397 12545
rect 5355 12496 5356 12536
rect 5396 12496 5397 12536
rect 5355 12487 5397 12496
rect 33867 12536 33909 12545
rect 33867 12496 33868 12536
rect 33908 12496 33909 12536
rect 33867 12487 33909 12496
rect 34243 12536 34301 12537
rect 34243 12496 34252 12536
rect 34292 12496 34301 12536
rect 34243 12495 34301 12496
rect 35107 12536 35165 12537
rect 35107 12496 35116 12536
rect 35156 12496 35165 12536
rect 35107 12495 35165 12496
rect 36747 12536 36789 12545
rect 36747 12496 36748 12536
rect 36788 12496 36789 12536
rect 36747 12487 36789 12496
rect 36843 12536 36885 12545
rect 36843 12496 36844 12536
rect 36884 12496 36885 12536
rect 36843 12487 36885 12496
rect 37123 12536 37181 12537
rect 37123 12496 37132 12536
rect 37172 12496 37181 12536
rect 37123 12495 37181 12496
rect 39051 12536 39093 12545
rect 39051 12496 39052 12536
rect 39092 12496 39093 12536
rect 39051 12487 39093 12496
rect 39427 12536 39485 12537
rect 39427 12496 39436 12536
rect 39476 12496 39485 12536
rect 39427 12495 39485 12496
rect 40291 12536 40349 12537
rect 40291 12496 40300 12536
rect 40340 12496 40349 12536
rect 40291 12495 40349 12496
rect 42211 12536 42269 12537
rect 42211 12496 42220 12536
rect 42260 12496 42269 12536
rect 42211 12495 42269 12496
rect 42411 12536 42453 12545
rect 42411 12496 42412 12536
rect 42452 12496 42453 12536
rect 42411 12487 42453 12496
rect 45483 12536 45525 12545
rect 45483 12496 45484 12536
rect 45524 12496 45525 12536
rect 45483 12487 45525 12496
rect 45859 12536 45917 12537
rect 45859 12496 45868 12536
rect 45908 12496 45917 12536
rect 45859 12495 45917 12496
rect 46723 12536 46781 12537
rect 46723 12496 46732 12536
rect 46772 12496 46781 12536
rect 46723 12495 46781 12496
rect 48163 12536 48221 12537
rect 48163 12496 48172 12536
rect 48212 12496 48221 12536
rect 48163 12495 48221 12496
rect 48459 12536 48501 12545
rect 48459 12496 48460 12536
rect 48500 12496 48501 12536
rect 48459 12487 48501 12496
rect 49035 12536 49077 12545
rect 49035 12496 49036 12536
rect 49076 12496 49077 12536
rect 49035 12487 49077 12496
rect 49227 12536 49269 12545
rect 49227 12496 49228 12536
rect 49268 12496 49269 12536
rect 49227 12487 49269 12496
rect 49315 12536 49373 12537
rect 49315 12496 49324 12536
rect 49364 12496 49373 12536
rect 49315 12495 49373 12496
rect 49507 12536 49565 12537
rect 49507 12496 49516 12536
rect 49556 12496 49565 12536
rect 49507 12495 49565 12496
rect 49611 12536 49653 12545
rect 49611 12496 49612 12536
rect 49652 12496 49653 12536
rect 49611 12487 49653 12496
rect 49707 12536 49749 12545
rect 49707 12496 49708 12536
rect 49748 12496 49749 12536
rect 49707 12487 49749 12496
rect 51619 12536 51677 12537
rect 51619 12496 51628 12536
rect 51668 12496 51677 12536
rect 51619 12495 51677 12496
rect 51819 12536 51861 12545
rect 51819 12496 51820 12536
rect 51860 12496 51861 12536
rect 51819 12487 51861 12496
rect 52011 12536 52053 12545
rect 52011 12496 52012 12536
rect 52052 12496 52053 12536
rect 52011 12487 52053 12496
rect 52387 12536 52445 12537
rect 52387 12496 52396 12536
rect 52436 12496 52445 12536
rect 52387 12495 52445 12496
rect 53251 12536 53309 12537
rect 53251 12496 53260 12536
rect 53300 12496 53309 12536
rect 53251 12495 53309 12496
rect 55267 12536 55325 12537
rect 55267 12496 55276 12536
rect 55316 12496 55325 12536
rect 55267 12495 55325 12496
rect 56131 12536 56189 12537
rect 56131 12496 56140 12536
rect 56180 12496 56189 12536
rect 56131 12495 56189 12496
rect 58243 12536 58301 12537
rect 58243 12496 58252 12536
rect 58292 12496 58301 12536
rect 58243 12495 58301 12496
rect 58443 12536 58485 12545
rect 58443 12496 58444 12536
rect 58484 12496 58485 12536
rect 58443 12487 58485 12496
rect 59307 12536 59349 12545
rect 59307 12496 59308 12536
rect 59348 12496 59349 12536
rect 59307 12487 59349 12496
rect 59491 12536 59549 12537
rect 59491 12496 59500 12536
rect 59540 12496 59549 12536
rect 59491 12495 59549 12496
rect 61323 12536 61365 12545
rect 61323 12496 61324 12536
rect 61364 12496 61365 12536
rect 61323 12487 61365 12496
rect 61515 12536 61557 12545
rect 61515 12496 61516 12536
rect 61556 12496 61557 12536
rect 61515 12487 61557 12496
rect 61603 12536 61661 12537
rect 61603 12496 61612 12536
rect 61652 12496 61661 12536
rect 61603 12495 61661 12496
rect 62091 12536 62133 12545
rect 62091 12496 62092 12536
rect 62132 12496 62133 12536
rect 62091 12487 62133 12496
rect 62283 12536 62325 12545
rect 62283 12496 62284 12536
rect 62324 12496 62325 12536
rect 62283 12487 62325 12496
rect 62371 12536 62429 12537
rect 62371 12496 62380 12536
rect 62420 12496 62429 12536
rect 62371 12495 62429 12496
rect 63051 12536 63093 12545
rect 63051 12496 63052 12536
rect 63092 12496 63093 12536
rect 63051 12487 63093 12496
rect 63243 12536 63285 12545
rect 63243 12496 63244 12536
rect 63284 12496 63285 12536
rect 63243 12487 63285 12496
rect 63331 12536 63389 12537
rect 63331 12496 63340 12536
rect 63380 12496 63389 12536
rect 63331 12495 63389 12496
rect 64387 12536 64445 12537
rect 64387 12496 64396 12536
rect 64436 12496 64445 12536
rect 64387 12495 64445 12496
rect 64587 12536 64629 12545
rect 64587 12496 64588 12536
rect 64628 12496 64629 12536
rect 64587 12487 64629 12496
rect 64779 12536 64821 12545
rect 64779 12496 64780 12536
rect 64820 12496 64821 12536
rect 64779 12487 64821 12496
rect 65155 12536 65213 12537
rect 65155 12496 65164 12536
rect 65204 12496 65213 12536
rect 65155 12495 65213 12496
rect 66019 12536 66077 12537
rect 66019 12496 66028 12536
rect 66068 12496 66077 12536
rect 66019 12495 66077 12496
rect 67371 12536 67413 12545
rect 67371 12496 67372 12536
rect 67412 12496 67413 12536
rect 67371 12487 67413 12496
rect 67747 12536 67805 12537
rect 67747 12496 67756 12536
rect 67796 12496 67805 12536
rect 67747 12495 67805 12496
rect 68611 12536 68669 12537
rect 68611 12496 68620 12536
rect 68660 12496 68669 12536
rect 68611 12495 68669 12496
rect 69955 12536 70013 12537
rect 69955 12496 69964 12536
rect 70004 12496 70013 12536
rect 69955 12495 70013 12496
rect 70059 12536 70101 12545
rect 70059 12496 70060 12536
rect 70100 12496 70101 12536
rect 70059 12487 70101 12496
rect 70251 12536 70293 12545
rect 70251 12496 70252 12536
rect 70292 12496 70293 12536
rect 70251 12487 70293 12496
rect 70443 12536 70485 12545
rect 70443 12496 70444 12536
rect 70484 12496 70485 12536
rect 70443 12487 70485 12496
rect 70819 12536 70877 12537
rect 70819 12496 70828 12536
rect 70868 12496 70877 12536
rect 70819 12495 70877 12496
rect 71683 12536 71741 12537
rect 71683 12496 71692 12536
rect 71732 12496 71741 12536
rect 71683 12495 71741 12496
rect 74283 12536 74325 12545
rect 74283 12496 74284 12536
rect 74324 12496 74325 12536
rect 74283 12487 74325 12496
rect 74475 12536 74517 12545
rect 74763 12538 74764 12578
rect 74804 12538 74805 12578
rect 76107 12580 76108 12620
rect 76148 12580 76149 12620
rect 76107 12571 76149 12580
rect 74475 12496 74476 12536
rect 74516 12496 74517 12536
rect 74475 12487 74517 12496
rect 74563 12536 74621 12537
rect 74563 12496 74572 12536
rect 74612 12496 74621 12536
rect 74763 12529 74805 12538
rect 74955 12536 74997 12545
rect 74563 12495 74621 12496
rect 74955 12496 74956 12536
rect 74996 12496 74997 12536
rect 74955 12487 74997 12496
rect 75043 12536 75101 12537
rect 75043 12496 75052 12536
rect 75092 12496 75101 12536
rect 75043 12495 75101 12496
rect 76003 12536 76061 12537
rect 76003 12496 76012 12536
rect 76052 12496 76061 12536
rect 76003 12495 76061 12496
rect 76203 12536 76245 12545
rect 76203 12496 76204 12536
rect 76244 12496 76245 12536
rect 76203 12487 76245 12496
rect 76875 12536 76917 12545
rect 76875 12496 76876 12536
rect 76916 12496 76917 12536
rect 76875 12487 76917 12496
rect 77251 12536 77309 12537
rect 77251 12496 77260 12536
rect 77300 12496 77309 12536
rect 77251 12495 77309 12496
rect 78115 12536 78173 12537
rect 78115 12496 78124 12536
rect 78164 12496 78173 12536
rect 78115 12495 78173 12496
rect 2187 12442 2229 12451
rect 36267 12452 36309 12461
rect 1699 12411 1757 12412
rect 36267 12412 36268 12452
rect 36308 12412 36309 12452
rect 36267 12403 36309 12412
rect 54411 12452 54453 12461
rect 54411 12412 54412 12452
rect 54452 12412 54453 12452
rect 54411 12403 54453 12412
rect 57859 12452 57917 12453
rect 57859 12412 57868 12452
rect 57908 12412 57917 12452
rect 57859 12411 57917 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 1131 12368 1173 12377
rect 1131 12328 1132 12368
rect 1172 12328 1173 12368
rect 1131 12319 1173 12328
rect 2379 12368 2421 12377
rect 2379 12328 2380 12368
rect 2420 12328 2421 12368
rect 2379 12319 2421 12328
rect 2859 12368 2901 12377
rect 2859 12328 2860 12368
rect 2900 12328 2901 12368
rect 2859 12319 2901 12328
rect 5931 12368 5973 12377
rect 5931 12328 5932 12368
rect 5972 12328 5973 12368
rect 5931 12319 5973 12328
rect 36451 12368 36509 12369
rect 36451 12328 36460 12368
rect 36500 12328 36509 12368
rect 36451 12327 36509 12328
rect 37419 12368 37461 12377
rect 37419 12328 37420 12368
rect 37460 12328 37461 12368
rect 37419 12319 37461 12328
rect 42795 12368 42837 12377
rect 42795 12328 42796 12368
rect 42836 12328 42837 12368
rect 42795 12319 42837 12328
rect 48835 12368 48893 12369
rect 48835 12328 48844 12368
rect 48884 12328 48893 12368
rect 48835 12327 48893 12328
rect 49899 12368 49941 12377
rect 49899 12328 49900 12368
rect 49940 12328 49941 12368
rect 49899 12319 49941 12328
rect 58347 12368 58389 12377
rect 58347 12328 58348 12368
rect 58388 12328 58389 12368
rect 58347 12319 58389 12328
rect 59787 12368 59829 12377
rect 59787 12328 59788 12368
rect 59828 12328 59829 12368
rect 59787 12319 59829 12328
rect 62091 12368 62133 12377
rect 62091 12328 62092 12368
rect 62132 12328 62133 12368
rect 62091 12319 62133 12328
rect 70251 12368 70293 12377
rect 70251 12328 70252 12368
rect 70292 12328 70293 12368
rect 70251 12319 70293 12328
rect 74763 12368 74805 12377
rect 74763 12328 74764 12368
rect 74804 12328 74805 12368
rect 74763 12319 74805 12328
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 42315 12284 42357 12293
rect 42315 12244 42316 12284
rect 42356 12244 42357 12284
rect 42315 12235 42357 12244
rect 51723 12284 51765 12293
rect 51723 12244 51724 12284
rect 51764 12244 51765 12284
rect 51723 12235 51765 12244
rect 58059 12284 58101 12293
rect 58059 12244 58060 12284
rect 58100 12244 58101 12284
rect 58059 12235 58101 12244
rect 59403 12284 59445 12293
rect 59403 12244 59404 12284
rect 59444 12244 59445 12284
rect 59403 12235 59445 12244
rect 63051 12284 63093 12293
rect 63051 12244 63052 12284
rect 63092 12244 63093 12284
rect 63051 12235 63093 12244
rect 64491 12284 64533 12293
rect 64491 12244 64492 12284
rect 64532 12244 64533 12284
rect 64491 12235 64533 12244
rect 69763 12284 69821 12285
rect 69763 12244 69772 12284
rect 69812 12244 69821 12284
rect 69763 12243 69821 12244
rect 79267 12284 79325 12285
rect 79267 12244 79276 12284
rect 79316 12244 79325 12284
rect 79267 12243 79325 12244
rect 576 12116 79584 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 75112 12116
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75480 12076 79584 12116
rect 576 12052 79584 12076
rect 34827 11948 34869 11957
rect 34827 11908 34828 11948
rect 34868 11908 34869 11948
rect 34827 11899 34869 11908
rect 36843 11948 36885 11957
rect 36843 11908 36844 11948
rect 36884 11908 36885 11948
rect 36843 11899 36885 11908
rect 39435 11948 39477 11957
rect 39435 11908 39436 11948
rect 39476 11908 39477 11948
rect 39435 11899 39477 11908
rect 44707 11948 44765 11949
rect 44707 11908 44716 11948
rect 44756 11908 44765 11948
rect 44707 11907 44765 11908
rect 46827 11948 46869 11957
rect 46827 11908 46828 11948
rect 46868 11908 46869 11948
rect 46827 11899 46869 11908
rect 48267 11948 48309 11957
rect 48267 11908 48268 11948
rect 48308 11908 48309 11948
rect 48267 11899 48309 11908
rect 61699 11948 61757 11949
rect 61699 11908 61708 11948
rect 61748 11908 61757 11948
rect 61699 11907 61757 11908
rect 64587 11948 64629 11957
rect 64587 11908 64588 11948
rect 64628 11908 64629 11948
rect 64587 11899 64629 11908
rect 69475 11948 69533 11949
rect 69475 11908 69484 11948
rect 69524 11908 69533 11948
rect 69475 11907 69533 11908
rect 70539 11948 70581 11957
rect 70539 11908 70540 11948
rect 70580 11908 70581 11948
rect 70539 11899 70581 11908
rect 74851 11948 74909 11949
rect 74851 11908 74860 11948
rect 74900 11908 74909 11948
rect 74851 11907 74909 11908
rect 76395 11948 76437 11957
rect 76395 11908 76396 11948
rect 76436 11908 76437 11948
rect 76395 11899 76437 11908
rect 1227 11864 1269 11873
rect 1227 11824 1228 11864
rect 1268 11824 1269 11864
rect 1227 11815 1269 11824
rect 1803 11864 1845 11873
rect 1803 11824 1804 11864
rect 1844 11824 1845 11864
rect 1803 11815 1845 11824
rect 4003 11864 4061 11865
rect 4003 11824 4012 11864
rect 4052 11824 4061 11864
rect 4003 11823 4061 11824
rect 34347 11864 34389 11873
rect 34347 11824 34348 11864
rect 34388 11824 34389 11864
rect 34347 11815 34389 11824
rect 38467 11864 38525 11865
rect 38467 11824 38476 11864
rect 38516 11824 38525 11864
rect 38467 11823 38525 11824
rect 42123 11864 42165 11873
rect 42123 11824 42124 11864
rect 42164 11824 42165 11864
rect 42123 11815 42165 11824
rect 44907 11864 44949 11873
rect 44907 11824 44908 11864
rect 44948 11824 44949 11864
rect 44907 11815 44949 11824
rect 45963 11864 46005 11873
rect 45963 11824 45964 11864
rect 46004 11824 46005 11864
rect 45963 11815 46005 11824
rect 49131 11864 49173 11873
rect 49131 11824 49132 11864
rect 49172 11824 49173 11864
rect 49131 11815 49173 11824
rect 49803 11864 49845 11873
rect 49803 11824 49804 11864
rect 49844 11824 49845 11864
rect 49803 11815 49845 11824
rect 51427 11864 51485 11865
rect 51427 11824 51436 11864
rect 51476 11824 51485 11864
rect 51427 11823 51485 11824
rect 52491 11864 52533 11873
rect 52491 11824 52492 11864
rect 52532 11824 52533 11864
rect 52491 11815 52533 11824
rect 55371 11864 55413 11873
rect 55371 11824 55372 11864
rect 55412 11824 55413 11864
rect 55371 11815 55413 11824
rect 56331 11864 56373 11873
rect 56331 11824 56332 11864
rect 56372 11824 56373 11864
rect 56331 11815 56373 11824
rect 57291 11864 57333 11873
rect 57291 11824 57292 11864
rect 57332 11824 57333 11864
rect 57291 11815 57333 11824
rect 62091 11864 62133 11873
rect 62091 11824 62092 11864
rect 62132 11824 62133 11864
rect 62091 11815 62133 11824
rect 64099 11864 64157 11865
rect 64099 11824 64108 11864
rect 64148 11824 64157 11864
rect 64099 11823 64157 11824
rect 65355 11864 65397 11873
rect 65355 11824 65356 11864
rect 65396 11824 65397 11864
rect 65355 11815 65397 11824
rect 67563 11864 67605 11873
rect 67563 11824 67564 11864
rect 67604 11824 67605 11864
rect 67563 11815 67605 11824
rect 76003 11864 76061 11865
rect 76003 11824 76012 11864
rect 76052 11824 76061 11864
rect 76003 11823 76061 11824
rect 77355 11864 77397 11873
rect 77355 11824 77356 11864
rect 77396 11824 77397 11864
rect 77355 11815 77397 11824
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 1411 11780 1469 11781
rect 1411 11740 1420 11780
rect 1460 11740 1469 11780
rect 1411 11739 1469 11740
rect 7371 11780 7413 11789
rect 7371 11740 7372 11780
rect 7412 11740 7413 11780
rect 7371 11731 7413 11740
rect 49603 11780 49661 11781
rect 49603 11740 49612 11780
rect 49652 11740 49661 11780
rect 49603 11739 49661 11740
rect 57475 11780 57533 11781
rect 57475 11740 57484 11780
rect 57524 11740 57533 11780
rect 57475 11739 57533 11740
rect 1995 11696 2037 11705
rect 1995 11656 1996 11696
rect 2036 11656 2037 11696
rect 1995 11647 2037 11656
rect 2091 11696 2133 11705
rect 2091 11656 2092 11696
rect 2132 11656 2133 11696
rect 2091 11647 2133 11656
rect 2187 11696 2229 11705
rect 2187 11656 2188 11696
rect 2228 11656 2229 11696
rect 2187 11647 2229 11656
rect 3331 11696 3389 11697
rect 3331 11656 3340 11696
rect 3380 11656 3389 11696
rect 3331 11655 3389 11656
rect 3627 11696 3669 11705
rect 3627 11656 3628 11696
rect 3668 11656 3669 11696
rect 3627 11647 3669 11656
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 4491 11696 4533 11705
rect 4491 11656 4492 11696
rect 4532 11656 4533 11696
rect 4491 11647 4533 11656
rect 4683 11696 4725 11705
rect 4683 11656 4684 11696
rect 4724 11656 4725 11696
rect 4683 11647 4725 11656
rect 4771 11696 4829 11697
rect 4771 11656 4780 11696
rect 4820 11656 4829 11696
rect 4771 11655 4829 11656
rect 4971 11696 5013 11705
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 5347 11696 5405 11697
rect 5347 11656 5356 11696
rect 5396 11656 5405 11696
rect 5347 11655 5405 11656
rect 6211 11696 6269 11697
rect 6211 11656 6220 11696
rect 6260 11656 6269 11696
rect 6211 11655 6269 11656
rect 34827 11696 34869 11705
rect 34827 11656 34828 11696
rect 34868 11656 34869 11696
rect 34827 11647 34869 11656
rect 35019 11696 35061 11705
rect 35019 11656 35020 11696
rect 35060 11656 35061 11696
rect 35019 11647 35061 11656
rect 35107 11696 35165 11697
rect 35107 11656 35116 11696
rect 35156 11656 35165 11696
rect 35107 11655 35165 11656
rect 35307 11696 35349 11705
rect 35307 11656 35308 11696
rect 35348 11656 35349 11696
rect 35307 11647 35349 11656
rect 35403 11696 35445 11705
rect 35403 11656 35404 11696
rect 35444 11656 35445 11696
rect 35403 11647 35445 11656
rect 35499 11696 35541 11705
rect 35499 11656 35500 11696
rect 35540 11656 35541 11696
rect 35499 11647 35541 11656
rect 35595 11696 35637 11705
rect 35595 11656 35596 11696
rect 35636 11656 35637 11696
rect 35595 11647 35637 11656
rect 36067 11696 36125 11697
rect 36067 11656 36076 11696
rect 36116 11656 36125 11696
rect 36067 11655 36125 11656
rect 36171 11696 36213 11705
rect 36171 11656 36172 11696
rect 36212 11656 36213 11696
rect 36171 11647 36213 11656
rect 36363 11696 36405 11705
rect 36363 11656 36364 11696
rect 36404 11656 36405 11696
rect 36363 11647 36405 11656
rect 36547 11696 36605 11697
rect 36547 11656 36556 11696
rect 36596 11656 36605 11696
rect 36547 11655 36605 11656
rect 36651 11696 36693 11705
rect 36651 11656 36652 11696
rect 36692 11656 36693 11696
rect 36651 11647 36693 11656
rect 36843 11696 36885 11705
rect 36843 11656 36844 11696
rect 36884 11656 36885 11696
rect 36843 11647 36885 11656
rect 38083 11696 38141 11697
rect 38083 11656 38092 11696
rect 38132 11656 38141 11696
rect 38083 11655 38141 11656
rect 38283 11696 38325 11705
rect 38283 11656 38284 11696
rect 38324 11656 38325 11696
rect 38283 11647 38325 11656
rect 38859 11696 38901 11705
rect 38859 11656 38860 11696
rect 38900 11656 38901 11696
rect 38859 11647 38901 11656
rect 39139 11696 39197 11697
rect 39139 11656 39148 11696
rect 39188 11656 39197 11696
rect 39139 11655 39197 11656
rect 39435 11696 39477 11705
rect 39435 11656 39436 11696
rect 39476 11656 39477 11696
rect 39435 11647 39477 11656
rect 39627 11696 39669 11705
rect 39627 11656 39628 11696
rect 39668 11656 39669 11696
rect 39627 11647 39669 11656
rect 39715 11696 39773 11697
rect 39715 11656 39724 11696
rect 39764 11656 39773 11696
rect 39715 11655 39773 11656
rect 41827 11696 41885 11697
rect 41827 11656 41836 11696
rect 41876 11656 41885 11696
rect 41827 11655 41885 11656
rect 41931 11696 41973 11705
rect 41931 11656 41932 11696
rect 41972 11656 41973 11696
rect 41931 11647 41973 11656
rect 42123 11696 42165 11705
rect 42123 11656 42124 11696
rect 42164 11656 42165 11696
rect 42123 11647 42165 11656
rect 42315 11696 42357 11705
rect 42315 11656 42316 11696
rect 42356 11656 42357 11696
rect 42315 11647 42357 11656
rect 42691 11696 42749 11697
rect 42691 11656 42700 11696
rect 42740 11656 42749 11696
rect 42691 11655 42749 11656
rect 43555 11696 43613 11697
rect 43555 11656 43564 11696
rect 43604 11656 43613 11696
rect 43555 11655 43613 11656
rect 46347 11696 46389 11705
rect 46347 11656 46348 11696
rect 46388 11656 46389 11696
rect 46347 11647 46389 11656
rect 46443 11696 46485 11705
rect 46443 11656 46444 11696
rect 46484 11656 46485 11696
rect 46443 11647 46485 11656
rect 46539 11696 46581 11705
rect 46539 11656 46540 11696
rect 46580 11656 46581 11696
rect 46539 11647 46581 11656
rect 46635 11696 46677 11705
rect 46635 11656 46636 11696
rect 46676 11656 46677 11696
rect 46635 11647 46677 11656
rect 46827 11696 46869 11705
rect 46827 11656 46828 11696
rect 46868 11656 46869 11696
rect 46827 11647 46869 11656
rect 47019 11696 47061 11705
rect 47019 11656 47020 11696
rect 47060 11656 47061 11696
rect 47019 11647 47061 11656
rect 47107 11696 47165 11697
rect 47107 11656 47116 11696
rect 47156 11656 47165 11696
rect 47107 11655 47165 11656
rect 48267 11696 48309 11705
rect 48267 11656 48268 11696
rect 48308 11656 48309 11696
rect 48267 11647 48309 11656
rect 48459 11696 48501 11705
rect 48459 11656 48460 11696
rect 48500 11656 48501 11696
rect 48459 11647 48501 11656
rect 48547 11696 48605 11697
rect 48547 11656 48556 11696
rect 48596 11656 48605 11696
rect 48547 11655 48605 11656
rect 49131 11696 49173 11705
rect 49131 11656 49132 11696
rect 49172 11656 49173 11696
rect 49131 11647 49173 11656
rect 49323 11696 49365 11705
rect 49323 11656 49324 11696
rect 49364 11656 49365 11696
rect 49323 11647 49365 11656
rect 49411 11696 49469 11697
rect 49411 11656 49420 11696
rect 49460 11656 49469 11696
rect 50283 11696 50325 11705
rect 49411 11655 49469 11656
rect 50187 11675 50229 11684
rect 50187 11635 50188 11675
rect 50228 11635 50229 11675
rect 50283 11656 50284 11696
rect 50324 11656 50325 11696
rect 50283 11647 50325 11656
rect 50379 11696 50421 11705
rect 50379 11656 50380 11696
rect 50420 11656 50421 11696
rect 50379 11647 50421 11656
rect 50755 11696 50813 11697
rect 50755 11656 50764 11696
rect 50804 11656 50813 11696
rect 50755 11655 50813 11656
rect 51051 11696 51093 11705
rect 51051 11656 51052 11696
rect 51092 11656 51093 11696
rect 51051 11647 51093 11656
rect 51619 11696 51677 11697
rect 51619 11656 51628 11696
rect 51668 11656 51677 11696
rect 51619 11655 51677 11656
rect 51723 11696 51765 11705
rect 51723 11656 51724 11696
rect 51764 11656 51765 11696
rect 51723 11647 51765 11656
rect 51915 11696 51957 11705
rect 51915 11656 51916 11696
rect 51956 11656 51957 11696
rect 51915 11647 51957 11656
rect 53731 11696 53789 11697
rect 53731 11656 53740 11696
rect 53780 11656 53789 11696
rect 53731 11655 53789 11656
rect 53931 11696 53973 11705
rect 53931 11656 53932 11696
rect 53972 11656 53973 11696
rect 53931 11647 53973 11656
rect 56523 11696 56565 11705
rect 56523 11656 56524 11696
rect 56564 11656 56565 11696
rect 56523 11647 56565 11656
rect 56619 11696 56661 11705
rect 56619 11656 56620 11696
rect 56660 11656 56661 11696
rect 56619 11647 56661 11656
rect 56715 11696 56757 11705
rect 56715 11656 56716 11696
rect 56756 11656 56757 11696
rect 56715 11647 56757 11656
rect 56811 11696 56853 11705
rect 56811 11656 56812 11696
rect 56852 11656 56853 11696
rect 56811 11647 56853 11656
rect 57675 11696 57717 11705
rect 57675 11656 57676 11696
rect 57716 11656 57717 11696
rect 57675 11647 57717 11656
rect 57867 11696 57909 11705
rect 57867 11656 57868 11696
rect 57908 11656 57909 11696
rect 57867 11647 57909 11656
rect 57955 11696 58013 11697
rect 57955 11656 57964 11696
rect 58004 11656 58013 11696
rect 57955 11655 58013 11656
rect 58251 11696 58293 11705
rect 58251 11656 58252 11696
rect 58292 11656 58293 11696
rect 58251 11647 58293 11656
rect 58347 11696 58389 11705
rect 58347 11656 58348 11696
rect 58388 11656 58389 11696
rect 58347 11647 58389 11656
rect 58443 11696 58485 11705
rect 58443 11656 58444 11696
rect 58484 11656 58485 11696
rect 58443 11647 58485 11656
rect 58827 11696 58869 11705
rect 58827 11656 58828 11696
rect 58868 11656 58869 11696
rect 58827 11647 58869 11656
rect 59019 11696 59061 11705
rect 59019 11656 59020 11696
rect 59060 11656 59061 11696
rect 59019 11647 59061 11656
rect 59107 11696 59165 11697
rect 59107 11656 59116 11696
rect 59156 11656 59165 11696
rect 59107 11655 59165 11656
rect 59683 11696 59741 11697
rect 59683 11656 59692 11696
rect 59732 11656 59741 11696
rect 59683 11655 59741 11656
rect 60547 11696 60605 11697
rect 60547 11656 60556 11696
rect 60596 11656 60605 11696
rect 62859 11696 62901 11705
rect 60547 11655 60605 11656
rect 62763 11675 62805 11684
rect 50187 11626 50229 11635
rect 62763 11635 62764 11675
rect 62804 11635 62805 11675
rect 62859 11656 62860 11696
rect 62900 11656 62901 11696
rect 62859 11647 62901 11656
rect 62955 11696 62997 11705
rect 62955 11656 62956 11696
rect 62996 11656 62997 11696
rect 62955 11647 62997 11656
rect 63051 11696 63093 11705
rect 63051 11656 63052 11696
rect 63092 11656 63093 11696
rect 63051 11647 63093 11656
rect 63427 11696 63485 11697
rect 63427 11656 63436 11696
rect 63476 11656 63485 11696
rect 63427 11655 63485 11656
rect 63723 11696 63765 11705
rect 63723 11656 63724 11696
rect 63764 11656 63765 11696
rect 63723 11647 63765 11656
rect 64291 11696 64349 11697
rect 64291 11656 64300 11696
rect 64340 11656 64349 11696
rect 64291 11655 64349 11656
rect 64395 11696 64437 11705
rect 64395 11656 64396 11696
rect 64436 11656 64437 11696
rect 64395 11647 64437 11656
rect 64587 11696 64629 11705
rect 64587 11656 64588 11696
rect 64628 11656 64629 11696
rect 64587 11647 64629 11656
rect 68907 11696 68949 11705
rect 68907 11656 68908 11696
rect 68948 11656 68949 11696
rect 68907 11647 68949 11656
rect 69099 11696 69141 11705
rect 69099 11656 69100 11696
rect 69140 11656 69141 11696
rect 69099 11647 69141 11656
rect 69187 11696 69245 11697
rect 69187 11656 69196 11696
rect 69236 11656 69245 11696
rect 69187 11655 69245 11656
rect 69867 11696 69909 11705
rect 69867 11656 69868 11696
rect 69908 11656 69909 11696
rect 69867 11647 69909 11656
rect 70147 11696 70205 11697
rect 70147 11656 70156 11696
rect 70196 11656 70205 11696
rect 70147 11655 70205 11656
rect 70435 11696 70493 11697
rect 70435 11656 70444 11696
rect 70484 11656 70493 11696
rect 70435 11655 70493 11656
rect 70635 11696 70677 11705
rect 70635 11656 70636 11696
rect 70676 11656 70677 11696
rect 70635 11647 70677 11656
rect 72835 11696 72893 11697
rect 72835 11656 72844 11696
rect 72884 11656 72893 11696
rect 72835 11655 72893 11656
rect 73699 11696 73757 11697
rect 73699 11656 73708 11696
rect 73748 11656 73757 11696
rect 73699 11655 73757 11656
rect 75331 11696 75389 11697
rect 75331 11656 75340 11696
rect 75380 11656 75389 11696
rect 75331 11655 75389 11656
rect 75627 11696 75669 11705
rect 75627 11656 75628 11696
rect 75668 11656 75669 11696
rect 75627 11647 75669 11656
rect 75723 11696 75765 11705
rect 75723 11656 75724 11696
rect 75764 11656 75765 11696
rect 75723 11647 75765 11656
rect 76395 11696 76437 11705
rect 76395 11656 76396 11696
rect 76436 11656 76437 11696
rect 76395 11647 76437 11656
rect 76587 11696 76629 11705
rect 76587 11656 76588 11696
rect 76628 11656 76629 11696
rect 76587 11647 76629 11656
rect 76675 11696 76733 11697
rect 76675 11656 76684 11696
rect 76724 11656 76733 11696
rect 76675 11655 76733 11656
rect 76867 11696 76925 11697
rect 76867 11656 76876 11696
rect 76916 11656 76925 11696
rect 76867 11655 76925 11656
rect 77067 11696 77109 11705
rect 77067 11656 77068 11696
rect 77108 11656 77109 11696
rect 77067 11647 77109 11656
rect 62763 11626 62805 11635
rect 4587 11612 4629 11621
rect 4587 11572 4588 11612
rect 4628 11572 4629 11612
rect 4587 11563 4629 11572
rect 38187 11612 38229 11621
rect 38187 11572 38188 11612
rect 38228 11572 38229 11612
rect 38187 11563 38229 11572
rect 38763 11612 38805 11621
rect 38763 11572 38764 11612
rect 38804 11572 38805 11612
rect 38763 11563 38805 11572
rect 51147 11612 51189 11621
rect 51147 11572 51148 11612
rect 51188 11572 51189 11612
rect 51147 11563 51189 11572
rect 51819 11612 51861 11621
rect 51819 11572 51820 11612
rect 51860 11572 51861 11612
rect 51819 11563 51861 11572
rect 53835 11612 53877 11621
rect 53835 11572 53836 11612
rect 53876 11572 53877 11612
rect 53835 11563 53877 11572
rect 58923 11612 58965 11621
rect 58923 11572 58924 11612
rect 58964 11572 58965 11612
rect 58923 11563 58965 11572
rect 59307 11612 59349 11621
rect 59307 11572 59308 11612
rect 59348 11572 59349 11612
rect 59307 11563 59349 11572
rect 63819 11612 63861 11621
rect 63819 11572 63820 11612
rect 63860 11572 63861 11612
rect 63819 11563 63861 11572
rect 69003 11612 69045 11621
rect 69003 11572 69004 11612
rect 69044 11572 69045 11612
rect 69003 11563 69045 11572
rect 69771 11612 69813 11621
rect 69771 11572 69772 11612
rect 69812 11572 69813 11612
rect 69771 11563 69813 11572
rect 72459 11612 72501 11621
rect 72459 11572 72460 11612
rect 72500 11572 72501 11612
rect 72459 11563 72501 11572
rect 76971 11612 77013 11621
rect 76971 11572 76972 11612
rect 77012 11572 77013 11612
rect 76971 11563 77013 11572
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 2275 11528 2333 11529
rect 2275 11488 2284 11528
rect 2324 11488 2333 11528
rect 2275 11487 2333 11488
rect 36259 11528 36317 11529
rect 36259 11488 36268 11528
rect 36308 11488 36317 11528
rect 36259 11487 36317 11488
rect 50467 11528 50525 11529
rect 50467 11488 50476 11528
rect 50516 11488 50525 11528
rect 50467 11487 50525 11488
rect 57763 11528 57821 11529
rect 57763 11488 57772 11528
rect 57812 11488 57821 11528
rect 57763 11487 57821 11488
rect 58147 11528 58205 11529
rect 58147 11488 58156 11528
rect 58196 11488 58205 11528
rect 58147 11487 58205 11488
rect 576 11360 79584 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 76352 11360
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76720 11320 79584 11360
rect 576 11296 79584 11320
rect 3907 11192 3965 11193
rect 3907 11152 3916 11192
rect 3956 11152 3965 11192
rect 3907 11151 3965 11152
rect 37803 11192 37845 11201
rect 37803 11152 37804 11192
rect 37844 11152 37845 11192
rect 37803 11143 37845 11152
rect 50467 11192 50525 11193
rect 50467 11152 50476 11192
rect 50516 11152 50525 11192
rect 50467 11151 50525 11152
rect 56227 11192 56285 11193
rect 56227 11152 56236 11192
rect 56276 11152 56285 11192
rect 56227 11151 56285 11152
rect 58819 11192 58877 11193
rect 58819 11152 58828 11192
rect 58868 11152 58877 11192
rect 58819 11151 58877 11152
rect 60931 11192 60989 11193
rect 60931 11152 60940 11192
rect 60980 11152 60989 11192
rect 60931 11151 60989 11152
rect 75235 11192 75293 11193
rect 75235 11152 75244 11192
rect 75284 11152 75293 11192
rect 75235 11151 75293 11152
rect 4971 11108 5013 11117
rect 4971 11068 4972 11108
rect 5012 11068 5013 11108
rect 4971 11059 5013 11068
rect 47019 11108 47061 11117
rect 47019 11068 47020 11108
rect 47060 11068 47061 11108
rect 47019 11059 47061 11068
rect 48075 11108 48117 11117
rect 48075 11068 48076 11108
rect 48116 11068 48117 11108
rect 48075 11059 48117 11068
rect 50859 11108 50901 11117
rect 50859 11068 50860 11108
rect 50900 11068 50901 11108
rect 50859 11059 50901 11068
rect 59307 11108 59349 11117
rect 59307 11068 59308 11108
rect 59348 11068 59349 11108
rect 59307 11059 59349 11068
rect 63339 11108 63381 11117
rect 63339 11068 63340 11108
rect 63380 11068 63381 11108
rect 63339 11059 63381 11068
rect 64011 11108 64053 11117
rect 64011 11068 64012 11108
rect 64052 11068 64053 11108
rect 64011 11059 64053 11068
rect 76203 11108 76245 11117
rect 76203 11068 76204 11108
rect 76244 11068 76245 11108
rect 76203 11059 76245 11068
rect 77058 11037 77100 11046
rect 1515 11024 1557 11033
rect 1515 10984 1516 11024
rect 1556 10984 1557 11024
rect 1515 10975 1557 10984
rect 1891 11024 1949 11025
rect 1891 10984 1900 11024
rect 1940 10984 1949 11024
rect 1891 10983 1949 10984
rect 2755 11024 2813 11025
rect 2755 10984 2764 11024
rect 2804 10984 2813 11024
rect 2755 10983 2813 10984
rect 4107 11024 4149 11033
rect 4107 10984 4108 11024
rect 4148 10984 4149 11024
rect 4107 10975 4149 10984
rect 4291 11024 4349 11025
rect 4291 10984 4300 11024
rect 4340 10984 4349 11024
rect 4291 10983 4349 10984
rect 4867 11024 4925 11025
rect 4867 10984 4876 11024
rect 4916 10984 4925 11024
rect 4867 10983 4925 10984
rect 5067 11024 5109 11033
rect 5067 10984 5068 11024
rect 5108 10984 5109 11024
rect 5067 10975 5109 10984
rect 36355 11024 36413 11025
rect 36355 10984 36364 11024
rect 36404 10984 36413 11024
rect 36355 10983 36413 10984
rect 36459 11024 36501 11033
rect 36459 10984 36460 11024
rect 36500 10984 36501 11024
rect 36459 10975 36501 10984
rect 36651 11024 36693 11033
rect 36651 10984 36652 11024
rect 36692 10984 36693 11024
rect 36651 10975 36693 10984
rect 36843 11024 36885 11033
rect 36843 10984 36844 11024
rect 36884 10984 36885 11024
rect 36843 10975 36885 10984
rect 36939 11024 36981 11033
rect 36939 10984 36940 11024
rect 36980 10984 36981 11024
rect 36939 10975 36981 10984
rect 37035 11024 37077 11033
rect 37035 10984 37036 11024
rect 37076 10984 37077 11024
rect 37035 10975 37077 10984
rect 37131 11024 37173 11033
rect 37131 10984 37132 11024
rect 37172 10984 37173 11024
rect 37131 10975 37173 10984
rect 39427 11024 39485 11025
rect 39427 10984 39436 11024
rect 39476 10984 39485 11024
rect 39427 10983 39485 10984
rect 41539 11024 41597 11025
rect 41539 10984 41548 11024
rect 41588 10984 41597 11024
rect 41539 10983 41597 10984
rect 41835 11024 41877 11033
rect 41835 10984 41836 11024
rect 41876 10984 41877 11024
rect 41835 10975 41877 10984
rect 41931 11024 41973 11033
rect 41931 10984 41932 11024
rect 41972 10984 41973 11024
rect 41931 10975 41973 10984
rect 42411 11024 42453 11033
rect 42411 10984 42412 11024
rect 42452 10984 42453 11024
rect 42411 10975 42453 10984
rect 42595 11024 42653 11025
rect 42595 10984 42604 11024
rect 42644 10984 42653 11024
rect 42595 10983 42653 10984
rect 43267 11024 43325 11025
rect 43267 10984 43276 11024
rect 43316 10984 43325 11024
rect 43267 10983 43325 10984
rect 43467 11024 43509 11033
rect 43467 10984 43468 11024
rect 43508 10984 43509 11024
rect 43467 10975 43509 10984
rect 43651 11024 43709 11025
rect 43651 10984 43660 11024
rect 43700 10984 43709 11024
rect 43651 10983 43709 10984
rect 43755 11024 43797 11033
rect 43755 10984 43756 11024
rect 43796 10984 43797 11024
rect 43755 10975 43797 10984
rect 43947 11024 43989 11033
rect 43947 10984 43948 11024
rect 43988 10984 43989 11024
rect 43947 10975 43989 10984
rect 44139 11024 44181 11033
rect 44139 10984 44140 11024
rect 44180 10984 44181 11024
rect 44139 10975 44181 10984
rect 44515 11024 44573 11025
rect 44515 10984 44524 11024
rect 44564 10984 44573 11024
rect 44515 10983 44573 10984
rect 45379 11024 45437 11025
rect 45379 10984 45388 11024
rect 45428 10984 45437 11024
rect 45379 10983 45437 10984
rect 46915 11024 46973 11025
rect 46915 10984 46924 11024
rect 46964 10984 46973 11024
rect 46915 10983 46973 10984
rect 47115 11024 47157 11033
rect 47115 10984 47116 11024
rect 47156 10984 47157 11024
rect 47115 10975 47157 10984
rect 48451 11024 48509 11025
rect 48451 10984 48460 11024
rect 48500 10984 48509 11024
rect 48451 10983 48509 10984
rect 49315 11024 49373 11025
rect 49315 10984 49324 11024
rect 49364 10984 49373 11024
rect 49315 10983 49373 10984
rect 50763 11024 50805 11033
rect 50763 10984 50764 11024
rect 50804 10984 50805 11024
rect 50763 10975 50805 10984
rect 50955 11024 50997 11033
rect 50955 10984 50956 11024
rect 50996 10984 50997 11024
rect 50955 10975 50997 10984
rect 51043 11024 51101 11025
rect 51043 10984 51052 11024
rect 51092 10984 51101 11024
rect 51043 10983 51101 10984
rect 51331 11024 51389 11025
rect 51331 10984 51340 11024
rect 51380 10984 51389 11024
rect 51331 10983 51389 10984
rect 51531 11024 51573 11033
rect 51531 10984 51532 11024
rect 51572 10984 51573 11024
rect 51531 10975 51573 10984
rect 53355 11024 53397 11033
rect 53355 10984 53356 11024
rect 53396 10984 53397 11024
rect 53355 10975 53397 10984
rect 53547 11024 53589 11033
rect 53547 10984 53548 11024
rect 53588 10984 53589 11024
rect 53547 10975 53589 10984
rect 53635 11024 53693 11025
rect 53635 10984 53644 11024
rect 53684 10984 53693 11024
rect 53635 10983 53693 10984
rect 53835 11024 53877 11033
rect 53835 10984 53836 11024
rect 53876 10984 53877 11024
rect 53835 10975 53877 10984
rect 54211 11024 54269 11025
rect 54211 10984 54220 11024
rect 54260 10984 54269 11024
rect 54211 10983 54269 10984
rect 55075 11024 55133 11025
rect 55075 10984 55084 11024
rect 55124 10984 55133 11024
rect 55075 10983 55133 10984
rect 56427 11024 56469 11033
rect 56427 10984 56428 11024
rect 56468 10984 56469 11024
rect 56427 10975 56469 10984
rect 56803 11024 56861 11025
rect 56803 10984 56812 11024
rect 56852 10984 56861 11024
rect 56803 10983 56861 10984
rect 57667 11024 57725 11025
rect 57667 10984 57676 11024
rect 57716 10984 57725 11024
rect 57667 10983 57725 10984
rect 59403 11024 59445 11033
rect 59403 10984 59404 11024
rect 59444 10984 59445 11024
rect 59403 10975 59445 10984
rect 59683 11024 59741 11025
rect 59683 10984 59692 11024
rect 59732 10984 59741 11024
rect 59683 10983 59741 10984
rect 62083 11024 62141 11025
rect 62083 10984 62092 11024
rect 62132 10984 62141 11024
rect 62083 10983 62141 10984
rect 62947 11024 63005 11025
rect 62947 10984 62956 11024
rect 62996 10984 63005 11024
rect 62947 10983 63005 10984
rect 63907 11024 63965 11025
rect 63907 10984 63916 11024
rect 63956 10984 63965 11024
rect 63907 10983 63965 10984
rect 64107 11024 64149 11033
rect 64107 10984 64108 11024
rect 64148 10984 64149 11024
rect 64107 10975 64149 10984
rect 64579 11024 64637 11025
rect 64579 10984 64588 11024
rect 64628 10984 64637 11024
rect 64579 10983 64637 10984
rect 64779 11024 64821 11033
rect 64779 10984 64780 11024
rect 64820 10984 64821 11024
rect 64779 10975 64821 10984
rect 64971 11024 65013 11033
rect 64971 10984 64972 11024
rect 65012 10984 65013 11024
rect 64971 10975 65013 10984
rect 65163 11024 65205 11033
rect 65163 10984 65164 11024
rect 65204 10984 65205 11024
rect 65163 10975 65205 10984
rect 65251 11024 65309 11025
rect 65251 10984 65260 11024
rect 65300 10984 65309 11024
rect 65251 10983 65309 10984
rect 69003 11024 69045 11033
rect 69003 10984 69004 11024
rect 69044 10984 69045 11024
rect 69003 10975 69045 10984
rect 69195 11024 69237 11033
rect 69195 10984 69196 11024
rect 69236 10984 69237 11024
rect 69195 10975 69237 10984
rect 69283 11024 69341 11025
rect 69283 10984 69292 11024
rect 69332 10984 69341 11024
rect 69283 10983 69341 10984
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 74763 11024 74805 11033
rect 74763 10984 74764 11024
rect 74804 10984 74805 11024
rect 74763 10975 74805 10984
rect 74859 11024 74901 11033
rect 74859 10984 74860 11024
rect 74900 10984 74901 11024
rect 74859 10975 74901 10984
rect 74955 11024 74997 11033
rect 74955 10984 74956 11024
rect 74996 10984 74997 11024
rect 74955 10975 74997 10984
rect 75147 11024 75189 11033
rect 75147 10984 75148 11024
rect 75188 10984 75189 11024
rect 75147 10975 75189 10984
rect 75339 11024 75381 11033
rect 75339 10984 75340 11024
rect 75380 10984 75381 11024
rect 75339 10975 75381 10984
rect 75427 11024 75485 11025
rect 75427 10984 75436 11024
rect 75476 10984 75485 11024
rect 75427 10983 75485 10984
rect 75627 11024 75669 11033
rect 75627 10984 75628 11024
rect 75668 10984 75669 11024
rect 75627 10975 75669 10984
rect 75819 11024 75861 11033
rect 75819 10984 75820 11024
rect 75860 10984 75861 11024
rect 75819 10975 75861 10984
rect 75907 11024 75965 11025
rect 75907 10984 75916 11024
rect 75956 10984 75965 11024
rect 75907 10983 75965 10984
rect 76107 11024 76149 11033
rect 76107 10984 76108 11024
rect 76148 10984 76149 11024
rect 76107 10975 76149 10984
rect 76291 11024 76349 11025
rect 76291 10984 76300 11024
rect 76340 10984 76349 11024
rect 77058 10997 77059 11037
rect 77099 10997 77100 11037
rect 77058 10988 77100 10997
rect 77251 11024 77309 11025
rect 76291 10983 76349 10984
rect 77251 10984 77260 11024
rect 77300 10984 77309 11024
rect 77251 10983 77309 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 1315 10940 1373 10941
rect 1315 10900 1324 10940
rect 1364 10900 1373 10940
rect 1315 10899 1373 10900
rect 51907 10940 51965 10941
rect 51907 10900 51916 10940
rect 51956 10900 51965 10940
rect 51907 10899 51965 10900
rect 68803 10940 68861 10941
rect 68803 10900 68812 10940
rect 68852 10900 68861 10940
rect 68803 10899 68861 10900
rect 69667 10940 69725 10941
rect 69667 10900 69676 10940
rect 69716 10900 69725 10940
rect 69667 10899 69725 10900
rect 70147 10940 70205 10941
rect 70147 10900 70156 10940
rect 70196 10900 70205 10940
rect 70147 10899 70205 10900
rect 70531 10940 70589 10941
rect 70531 10900 70540 10940
rect 70580 10900 70589 10940
rect 70531 10899 70589 10900
rect 71107 10940 71165 10941
rect 71107 10900 71116 10940
rect 71156 10900 71165 10940
rect 71107 10899 71165 10900
rect 76483 10940 76541 10941
rect 76483 10900 76492 10940
rect 76532 10900 76541 10940
rect 76483 10899 76541 10900
rect 1131 10856 1173 10865
rect 1131 10816 1132 10856
rect 1172 10816 1173 10856
rect 1131 10807 1173 10816
rect 36171 10856 36213 10865
rect 36171 10816 36172 10856
rect 36212 10816 36213 10856
rect 36171 10807 36213 10816
rect 39819 10856 39861 10865
rect 39819 10816 39820 10856
rect 39860 10816 39861 10856
rect 39819 10807 39861 10816
rect 42211 10856 42269 10857
rect 42211 10816 42220 10856
rect 42260 10816 42269 10856
rect 42211 10815 42269 10816
rect 43371 10856 43413 10865
rect 43371 10816 43372 10856
rect 43412 10816 43413 10856
rect 43371 10807 43413 10816
rect 43947 10856 43989 10865
rect 43947 10816 43948 10856
rect 43988 10816 43989 10856
rect 43947 10807 43989 10816
rect 46531 10856 46589 10857
rect 46531 10816 46540 10856
rect 46580 10816 46589 10856
rect 46531 10815 46589 10816
rect 47883 10856 47925 10865
rect 47883 10816 47884 10856
rect 47924 10816 47925 10856
rect 47883 10807 47925 10816
rect 51435 10856 51477 10865
rect 51435 10816 51436 10856
rect 51476 10816 51477 10856
rect 51435 10807 51477 10816
rect 65835 10856 65877 10865
rect 65835 10816 65836 10856
rect 65876 10816 65877 10856
rect 65835 10807 65877 10816
rect 71307 10856 71349 10865
rect 71307 10816 71308 10856
rect 71348 10816 71349 10856
rect 71307 10807 71349 10816
rect 72939 10856 72981 10865
rect 72939 10816 72940 10856
rect 72980 10816 72981 10856
rect 72939 10807 72981 10816
rect 75627 10856 75669 10865
rect 75627 10816 75628 10856
rect 75668 10816 75669 10856
rect 75627 10807 75669 10816
rect 77643 10856 77685 10865
rect 77643 10816 77644 10856
rect 77684 10816 77685 10856
rect 77643 10807 77685 10816
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 4203 10772 4245 10781
rect 4203 10732 4204 10772
rect 4244 10732 4245 10772
rect 4203 10723 4245 10732
rect 36651 10772 36693 10781
rect 36651 10732 36652 10772
rect 36692 10732 36693 10772
rect 36651 10723 36693 10732
rect 42507 10772 42549 10781
rect 42507 10732 42508 10772
rect 42548 10732 42549 10772
rect 42507 10723 42549 10732
rect 51723 10772 51765 10781
rect 51723 10732 51724 10772
rect 51764 10732 51765 10772
rect 51723 10723 51765 10732
rect 53355 10772 53397 10781
rect 53355 10732 53356 10772
rect 53396 10732 53397 10772
rect 53355 10723 53397 10732
rect 59011 10772 59069 10773
rect 59011 10732 59020 10772
rect 59060 10732 59069 10772
rect 59011 10731 59069 10732
rect 64683 10772 64725 10781
rect 64683 10732 64684 10772
rect 64724 10732 64725 10772
rect 64683 10723 64725 10732
rect 64971 10772 65013 10781
rect 64971 10732 64972 10772
rect 65012 10732 65013 10772
rect 64971 10723 65013 10732
rect 68619 10772 68661 10781
rect 68619 10732 68620 10772
rect 68660 10732 68661 10772
rect 68619 10723 68661 10732
rect 69003 10772 69045 10781
rect 69003 10732 69004 10772
rect 69044 10732 69045 10772
rect 69003 10723 69045 10732
rect 69483 10772 69525 10781
rect 69483 10732 69484 10772
rect 69524 10732 69525 10772
rect 69483 10723 69525 10732
rect 69963 10772 70005 10781
rect 69963 10732 69964 10772
rect 70004 10732 70005 10772
rect 69963 10723 70005 10732
rect 70731 10772 70773 10781
rect 70731 10732 70732 10772
rect 70772 10732 70773 10772
rect 70731 10723 70773 10732
rect 70923 10772 70965 10781
rect 70923 10732 70924 10772
rect 70964 10732 70965 10772
rect 70923 10723 70965 10732
rect 76683 10772 76725 10781
rect 76683 10732 76684 10772
rect 76724 10732 76725 10772
rect 76683 10723 76725 10732
rect 77163 10772 77205 10781
rect 77163 10732 77164 10772
rect 77204 10732 77205 10772
rect 77163 10723 77205 10732
rect 576 10604 79584 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 75112 10604
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75480 10564 79584 10604
rect 576 10540 79584 10564
rect 38755 10436 38813 10437
rect 38755 10396 38764 10436
rect 38804 10396 38813 10436
rect 38755 10395 38813 10396
rect 41731 10436 41789 10437
rect 41731 10396 41740 10436
rect 41780 10396 41789 10436
rect 41731 10395 41789 10396
rect 49123 10436 49181 10437
rect 49123 10396 49132 10436
rect 49172 10396 49181 10436
rect 49123 10395 49181 10396
rect 58059 10436 58101 10445
rect 58059 10396 58060 10436
rect 58100 10396 58101 10436
rect 58059 10387 58101 10396
rect 63435 10436 63477 10445
rect 63435 10396 63436 10436
rect 63476 10396 63477 10436
rect 63435 10387 63477 10396
rect 64963 10436 65021 10437
rect 64963 10396 64972 10436
rect 65012 10396 65021 10436
rect 64963 10395 65021 10396
rect 67651 10436 67709 10437
rect 67651 10396 67660 10436
rect 67700 10396 67709 10436
rect 67651 10395 67709 10396
rect 72835 10436 72893 10437
rect 72835 10396 72844 10436
rect 72884 10396 72893 10436
rect 72835 10395 72893 10396
rect 75811 10436 75869 10437
rect 75811 10396 75820 10436
rect 75860 10396 75869 10436
rect 75811 10395 75869 10396
rect 76867 10436 76925 10437
rect 76867 10396 76876 10436
rect 76916 10396 76925 10436
rect 76867 10395 76925 10396
rect 1515 10352 1557 10361
rect 1515 10312 1516 10352
rect 1556 10312 1557 10352
rect 1515 10303 1557 10312
rect 2187 10352 2229 10361
rect 2187 10312 2188 10352
rect 2228 10312 2229 10352
rect 2187 10303 2229 10312
rect 2667 10352 2709 10361
rect 2667 10312 2668 10352
rect 2708 10312 2709 10352
rect 2667 10303 2709 10312
rect 3147 10352 3189 10361
rect 3147 10312 3148 10352
rect 3188 10312 3189 10352
rect 3147 10303 3189 10312
rect 5259 10352 5301 10361
rect 5259 10312 5260 10352
rect 5300 10312 5301 10352
rect 5259 10303 5301 10312
rect 44131 10352 44189 10353
rect 44131 10312 44140 10352
rect 44180 10312 44189 10352
rect 44131 10311 44189 10312
rect 53347 10352 53405 10353
rect 53347 10312 53356 10352
rect 53396 10312 53405 10352
rect 53347 10311 53405 10312
rect 54315 10352 54357 10361
rect 54315 10312 54316 10352
rect 54356 10312 54357 10352
rect 54315 10303 54357 10312
rect 57579 10352 57621 10361
rect 57579 10312 57580 10352
rect 57620 10312 57621 10352
rect 57579 10303 57621 10312
rect 58731 10352 58773 10361
rect 58731 10312 58732 10352
rect 58772 10312 58773 10352
rect 58731 10303 58773 10312
rect 60267 10352 60309 10361
rect 60267 10312 60268 10352
rect 60308 10312 60309 10352
rect 60267 10303 60309 10312
rect 62379 10352 62421 10361
rect 62379 10312 62380 10352
rect 62420 10312 62421 10352
rect 62379 10303 62421 10312
rect 67851 10352 67893 10361
rect 67851 10312 67852 10352
rect 67892 10312 67893 10352
rect 67851 10303 67893 10312
rect 69955 10352 70013 10353
rect 69955 10312 69964 10352
rect 70004 10312 70013 10352
rect 69955 10311 70013 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 1699 10268 1757 10269
rect 1699 10228 1708 10268
rect 1748 10228 1757 10268
rect 1699 10227 1757 10228
rect 3331 10268 3389 10269
rect 3331 10228 3340 10268
rect 3380 10228 3389 10268
rect 3331 10227 3389 10228
rect 42115 10268 42173 10269
rect 42115 10228 42124 10268
rect 42164 10228 42173 10268
rect 42115 10227 42173 10228
rect 57379 10268 57437 10269
rect 57379 10228 57388 10268
rect 57428 10228 57437 10268
rect 57379 10227 57437 10228
rect 58915 10268 58973 10269
rect 58915 10228 58924 10268
rect 58964 10228 58973 10268
rect 58915 10227 58973 10228
rect 59491 10268 59549 10269
rect 59491 10228 59500 10268
rect 59540 10228 59549 10268
rect 59491 10227 59549 10228
rect 60067 10268 60125 10269
rect 60067 10228 60076 10268
rect 60116 10228 60125 10268
rect 60067 10227 60125 10228
rect 79467 10268 79509 10277
rect 79467 10228 79468 10268
rect 79508 10228 79509 10268
rect 79467 10219 79509 10228
rect 2187 10184 2229 10193
rect 2187 10144 2188 10184
rect 2228 10144 2229 10184
rect 2187 10135 2229 10144
rect 2379 10184 2421 10193
rect 2379 10144 2380 10184
rect 2420 10144 2421 10184
rect 2379 10135 2421 10144
rect 2467 10184 2525 10185
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 2467 10143 2525 10144
rect 2667 10184 2709 10193
rect 2667 10144 2668 10184
rect 2708 10144 2709 10184
rect 2947 10184 3005 10185
rect 2667 10135 2709 10144
rect 2859 10142 2901 10151
rect 2947 10144 2956 10184
rect 2996 10144 3005 10184
rect 2947 10143 3005 10144
rect 36363 10184 36405 10193
rect 36363 10144 36364 10184
rect 36404 10144 36405 10184
rect 2859 10102 2860 10142
rect 2900 10102 2901 10142
rect 36363 10135 36405 10144
rect 36739 10184 36797 10185
rect 36739 10144 36748 10184
rect 36788 10144 36797 10184
rect 36739 10143 36797 10144
rect 37603 10184 37661 10185
rect 37603 10144 37612 10184
rect 37652 10144 37661 10184
rect 37603 10143 37661 10144
rect 38947 10184 39005 10185
rect 38947 10144 38956 10184
rect 38996 10144 39005 10184
rect 38947 10143 39005 10144
rect 39147 10184 39189 10193
rect 39147 10144 39148 10184
rect 39188 10144 39189 10184
rect 39147 10135 39189 10144
rect 39715 10184 39773 10185
rect 39715 10144 39724 10184
rect 39764 10144 39773 10184
rect 39715 10143 39773 10144
rect 40579 10184 40637 10185
rect 40579 10144 40588 10184
rect 40628 10144 40637 10184
rect 40579 10143 40637 10144
rect 43459 10184 43517 10185
rect 43459 10144 43468 10184
rect 43508 10144 43517 10184
rect 43459 10143 43517 10144
rect 43755 10184 43797 10193
rect 43755 10144 43756 10184
rect 43796 10144 43797 10184
rect 43755 10135 43797 10144
rect 44331 10184 44373 10193
rect 44331 10144 44332 10184
rect 44372 10144 44373 10184
rect 44331 10135 44373 10144
rect 44515 10184 44573 10185
rect 44515 10144 44524 10184
rect 44564 10144 44573 10184
rect 44515 10143 44573 10144
rect 46251 10184 46293 10193
rect 46251 10144 46252 10184
rect 46292 10144 46293 10184
rect 46251 10135 46293 10144
rect 46443 10184 46485 10193
rect 46443 10144 46444 10184
rect 46484 10144 46485 10184
rect 46443 10135 46485 10144
rect 46531 10184 46589 10185
rect 46531 10144 46540 10184
rect 46580 10144 46589 10184
rect 46531 10143 46589 10144
rect 47107 10184 47165 10185
rect 47107 10144 47116 10184
rect 47156 10144 47165 10184
rect 47107 10143 47165 10144
rect 47971 10184 48029 10185
rect 47971 10144 47980 10184
rect 48020 10144 48029 10184
rect 47971 10143 48029 10144
rect 50275 10184 50333 10185
rect 50275 10144 50284 10184
rect 50324 10144 50333 10184
rect 50275 10143 50333 10144
rect 51139 10184 51197 10185
rect 51139 10144 51148 10184
rect 51188 10144 51197 10184
rect 51139 10143 51197 10144
rect 52675 10184 52733 10185
rect 52675 10144 52684 10184
rect 52724 10144 52733 10184
rect 52675 10143 52733 10144
rect 52971 10184 53013 10193
rect 52971 10144 52972 10184
rect 53012 10144 53013 10184
rect 52971 10135 53013 10144
rect 53547 10184 53589 10193
rect 53547 10144 53548 10184
rect 53588 10144 53589 10184
rect 53547 10135 53589 10144
rect 53731 10184 53789 10185
rect 53731 10144 53740 10184
rect 53780 10144 53789 10184
rect 53731 10143 53789 10144
rect 57763 10184 57821 10185
rect 57763 10144 57772 10184
rect 57812 10144 57821 10184
rect 57763 10143 57821 10144
rect 57867 10184 57909 10193
rect 57867 10144 57868 10184
rect 57908 10144 57909 10184
rect 57867 10135 57909 10144
rect 58059 10184 58101 10193
rect 58059 10144 58060 10184
rect 58100 10144 58101 10184
rect 58059 10135 58101 10144
rect 58251 10184 58293 10193
rect 58251 10144 58252 10184
rect 58292 10144 58293 10184
rect 58251 10135 58293 10144
rect 58443 10184 58485 10193
rect 58443 10144 58444 10184
rect 58484 10144 58485 10184
rect 58443 10135 58485 10144
rect 58531 10184 58589 10185
rect 58531 10144 58540 10184
rect 58580 10144 58589 10184
rect 58531 10143 58589 10144
rect 59115 10184 59157 10193
rect 59115 10144 59116 10184
rect 59156 10144 59157 10184
rect 59115 10135 59157 10144
rect 59299 10184 59357 10185
rect 59299 10144 59308 10184
rect 59348 10144 59357 10184
rect 59299 10143 59357 10144
rect 63435 10184 63477 10193
rect 63435 10144 63436 10184
rect 63476 10144 63477 10184
rect 63435 10135 63477 10144
rect 63627 10184 63669 10193
rect 63627 10144 63628 10184
rect 63668 10144 63669 10184
rect 63627 10135 63669 10144
rect 63715 10184 63773 10185
rect 63715 10144 63724 10184
rect 63764 10144 63773 10184
rect 63715 10143 63773 10144
rect 64291 10184 64349 10185
rect 64291 10144 64300 10184
rect 64340 10144 64349 10184
rect 64291 10143 64349 10144
rect 64587 10184 64629 10193
rect 64587 10144 64588 10184
rect 64628 10144 64629 10184
rect 64587 10135 64629 10144
rect 65259 10184 65301 10193
rect 65259 10144 65260 10184
rect 65300 10144 65301 10184
rect 65259 10135 65301 10144
rect 65635 10184 65693 10185
rect 65635 10144 65644 10184
rect 65684 10144 65693 10184
rect 65635 10143 65693 10144
rect 66499 10184 66557 10185
rect 66499 10144 66508 10184
rect 66548 10144 66557 10184
rect 66499 10143 66557 10144
rect 68235 10184 68277 10193
rect 68235 10144 68236 10184
rect 68276 10144 68277 10184
rect 68235 10135 68277 10144
rect 68331 10184 68373 10193
rect 68331 10144 68332 10184
rect 68372 10144 68373 10184
rect 68331 10135 68373 10144
rect 68427 10184 68469 10193
rect 68427 10144 68428 10184
rect 68468 10144 68469 10184
rect 68427 10135 68469 10144
rect 68523 10184 68565 10193
rect 68523 10144 68524 10184
rect 68564 10144 68565 10184
rect 68523 10135 68565 10144
rect 68715 10184 68757 10193
rect 68715 10144 68716 10184
rect 68756 10144 68757 10184
rect 68715 10135 68757 10144
rect 68907 10184 68949 10193
rect 68907 10144 68908 10184
rect 68948 10144 68949 10184
rect 68907 10135 68949 10144
rect 68995 10184 69053 10185
rect 68995 10144 69004 10184
rect 69044 10144 69053 10184
rect 68995 10143 69053 10144
rect 69283 10184 69341 10185
rect 69283 10144 69292 10184
rect 69332 10144 69341 10184
rect 69283 10143 69341 10144
rect 69579 10184 69621 10193
rect 69579 10144 69580 10184
rect 69620 10144 69621 10184
rect 69579 10135 69621 10144
rect 69675 10184 69717 10193
rect 69675 10144 69676 10184
rect 69716 10144 69717 10184
rect 69675 10135 69717 10144
rect 70819 10184 70877 10185
rect 70819 10144 70828 10184
rect 70868 10144 70877 10184
rect 70819 10143 70877 10144
rect 71683 10184 71741 10185
rect 71683 10144 71692 10184
rect 71732 10144 71741 10184
rect 71683 10143 71741 10144
rect 73795 10184 73853 10185
rect 73795 10144 73804 10184
rect 73844 10144 73853 10184
rect 73795 10143 73853 10144
rect 74659 10184 74717 10185
rect 74659 10144 74668 10184
rect 74708 10144 74717 10184
rect 74659 10143 74717 10144
rect 76195 10184 76253 10185
rect 76195 10144 76204 10184
rect 76244 10144 76253 10184
rect 76195 10143 76253 10144
rect 76491 10184 76533 10193
rect 76491 10144 76492 10184
rect 76532 10144 76533 10184
rect 76491 10135 76533 10144
rect 76587 10184 76629 10193
rect 76587 10144 76588 10184
rect 76628 10144 76629 10184
rect 76587 10135 76629 10144
rect 77443 10184 77501 10185
rect 77443 10144 77452 10184
rect 77492 10144 77501 10184
rect 77443 10143 77501 10144
rect 78307 10184 78365 10185
rect 78307 10144 78316 10184
rect 78356 10144 78365 10184
rect 78307 10143 78365 10144
rect 2859 10093 2901 10102
rect 39051 10100 39093 10109
rect 39051 10060 39052 10100
rect 39092 10060 39093 10100
rect 39051 10051 39093 10060
rect 39339 10100 39381 10109
rect 39339 10060 39340 10100
rect 39380 10060 39381 10100
rect 39339 10051 39381 10060
rect 43851 10100 43893 10109
rect 43851 10060 43852 10100
rect 43892 10060 43893 10100
rect 43851 10051 43893 10060
rect 44427 10100 44469 10109
rect 44427 10060 44428 10100
rect 44468 10060 44469 10100
rect 44427 10051 44469 10060
rect 46347 10100 46389 10109
rect 46347 10060 46348 10100
rect 46388 10060 46389 10100
rect 46347 10051 46389 10060
rect 46731 10100 46773 10109
rect 46731 10060 46732 10100
rect 46772 10060 46773 10100
rect 46731 10051 46773 10060
rect 49899 10100 49941 10109
rect 49899 10060 49900 10100
rect 49940 10060 49941 10100
rect 49899 10051 49941 10060
rect 53067 10100 53109 10109
rect 53067 10060 53068 10100
rect 53108 10060 53109 10100
rect 53067 10051 53109 10060
rect 53643 10100 53685 10109
rect 53643 10060 53644 10100
rect 53684 10060 53685 10100
rect 53643 10051 53685 10060
rect 59211 10100 59253 10109
rect 59211 10060 59212 10100
rect 59252 10060 59253 10100
rect 59211 10051 59253 10060
rect 64683 10100 64725 10109
rect 64683 10060 64684 10100
rect 64724 10060 64725 10100
rect 64683 10051 64725 10060
rect 68811 10100 68853 10109
rect 68811 10060 68812 10100
rect 68852 10060 68853 10100
rect 68811 10051 68853 10060
rect 70443 10100 70485 10109
rect 70443 10060 70444 10100
rect 70484 10060 70485 10100
rect 70443 10051 70485 10060
rect 73419 10100 73461 10109
rect 73419 10060 73420 10100
rect 73460 10060 73461 10100
rect 73419 10051 73461 10060
rect 77067 10100 77109 10109
rect 77067 10060 77068 10100
rect 77108 10060 77109 10100
rect 77067 10051 77109 10060
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 42315 10016 42357 10025
rect 42315 9976 42316 10016
rect 42356 9976 42357 10016
rect 42315 9967 42357 9976
rect 52291 10016 52349 10017
rect 52291 9976 52300 10016
rect 52340 9976 52349 10016
rect 52291 9975 52349 9976
rect 58339 10016 58397 10017
rect 58339 9976 58348 10016
rect 58388 9976 58397 10016
rect 58339 9975 58397 9976
rect 59691 10016 59733 10025
rect 59691 9976 59692 10016
rect 59732 9976 59733 10016
rect 59691 9967 59733 9976
rect 59883 10016 59925 10025
rect 59883 9976 59884 10016
rect 59924 9976 59925 10016
rect 59883 9967 59925 9976
rect 75811 10016 75869 10017
rect 75811 9976 75820 10016
rect 75860 9976 75869 10016
rect 75811 9975 75869 9976
rect 576 9848 79584 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 76352 9848
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76720 9808 79584 9848
rect 576 9784 79584 9808
rect 1515 9680 1557 9689
rect 1515 9640 1516 9680
rect 1556 9640 1557 9680
rect 1515 9631 1557 9640
rect 7171 9680 7229 9681
rect 7171 9640 7180 9680
rect 7220 9640 7229 9680
rect 7171 9639 7229 9640
rect 40099 9680 40157 9681
rect 40099 9640 40108 9680
rect 40148 9640 40157 9680
rect 40099 9639 40157 9640
rect 52683 9680 52725 9689
rect 52683 9640 52684 9680
rect 52724 9640 52725 9680
rect 52683 9631 52725 9640
rect 53059 9680 53117 9681
rect 53059 9640 53068 9680
rect 53108 9640 53117 9680
rect 53059 9639 53117 9640
rect 61987 9680 62045 9681
rect 61987 9640 61996 9680
rect 62036 9640 62045 9680
rect 61987 9639 62045 9640
rect 64579 9680 64637 9681
rect 64579 9640 64588 9680
rect 64628 9640 64637 9680
rect 64579 9639 64637 9640
rect 69283 9680 69341 9681
rect 69283 9640 69292 9680
rect 69332 9640 69341 9680
rect 69283 9639 69341 9640
rect 69675 9680 69717 9689
rect 69675 9640 69676 9680
rect 69716 9640 69717 9680
rect 69675 9631 69717 9640
rect 75523 9680 75581 9681
rect 75523 9640 75532 9680
rect 75572 9640 75581 9680
rect 75523 9639 75581 9640
rect 77155 9680 77213 9681
rect 77155 9640 77164 9680
rect 77204 9640 77213 9680
rect 77155 9639 77213 9640
rect 4491 9596 4533 9605
rect 4491 9556 4492 9596
rect 4532 9556 4533 9596
rect 4491 9547 4533 9556
rect 4779 9596 4821 9605
rect 4779 9556 4780 9596
rect 4820 9556 4821 9596
rect 4779 9547 4821 9556
rect 62187 9596 62229 9605
rect 62187 9556 62188 9596
rect 62228 9556 62229 9596
rect 62187 9547 62229 9556
rect 64875 9596 64917 9605
rect 64875 9556 64876 9596
rect 64916 9556 64917 9596
rect 64875 9547 64917 9556
rect 65355 9596 65397 9605
rect 65355 9556 65356 9596
rect 65396 9556 65397 9596
rect 65355 9547 65397 9556
rect 66891 9596 66933 9605
rect 66891 9556 66892 9596
rect 66932 9556 66933 9596
rect 66891 9547 66933 9556
rect 75723 9533 75765 9542
rect 2851 9527 2909 9528
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2091 9512 2133 9521
rect 2091 9472 2092 9512
rect 2132 9472 2133 9512
rect 2091 9463 2133 9472
rect 2187 9512 2229 9521
rect 2187 9472 2188 9512
rect 2228 9472 2229 9512
rect 2187 9463 2229 9472
rect 2283 9512 2325 9521
rect 2283 9472 2284 9512
rect 2324 9472 2325 9512
rect 2851 9487 2860 9527
rect 2900 9487 2909 9527
rect 2851 9486 2909 9487
rect 3147 9512 3189 9521
rect 2283 9463 2325 9472
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 3907 9512 3965 9513
rect 3907 9472 3916 9512
rect 3956 9472 3965 9512
rect 3907 9471 3965 9472
rect 4291 9512 4349 9513
rect 4291 9472 4300 9512
rect 4340 9472 4349 9512
rect 4291 9471 4349 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 5155 9512 5213 9513
rect 5155 9472 5164 9512
rect 5204 9472 5213 9512
rect 5155 9471 5213 9472
rect 6019 9512 6077 9513
rect 6019 9472 6028 9512
rect 6068 9472 6077 9512
rect 6019 9471 6077 9472
rect 39139 9512 39197 9513
rect 39139 9472 39148 9512
rect 39188 9472 39197 9512
rect 39139 9471 39197 9472
rect 39243 9512 39285 9521
rect 39243 9472 39244 9512
rect 39284 9472 39285 9512
rect 39243 9463 39285 9472
rect 39435 9512 39477 9521
rect 39435 9472 39436 9512
rect 39476 9472 39477 9512
rect 39435 9463 39477 9472
rect 39907 9512 39965 9513
rect 39907 9472 39916 9512
rect 39956 9472 39965 9512
rect 39907 9471 39965 9472
rect 40011 9512 40053 9521
rect 40011 9472 40012 9512
rect 40052 9472 40053 9512
rect 40011 9463 40053 9472
rect 40203 9512 40245 9521
rect 40203 9472 40204 9512
rect 40244 9472 40245 9512
rect 40203 9463 40245 9472
rect 40587 9512 40629 9521
rect 40587 9472 40588 9512
rect 40628 9472 40629 9512
rect 40587 9463 40629 9472
rect 40683 9512 40725 9521
rect 40683 9472 40684 9512
rect 40724 9472 40725 9512
rect 40683 9463 40725 9472
rect 40779 9512 40821 9521
rect 40779 9472 40780 9512
rect 40820 9472 40821 9512
rect 40779 9463 40821 9472
rect 40875 9512 40917 9521
rect 40875 9472 40876 9512
rect 40916 9472 40917 9512
rect 40875 9463 40917 9472
rect 41635 9512 41693 9513
rect 41635 9472 41644 9512
rect 41684 9472 41693 9512
rect 41635 9471 41693 9472
rect 41739 9512 41781 9521
rect 41739 9472 41740 9512
rect 41780 9472 41781 9512
rect 41739 9463 41781 9472
rect 41931 9512 41973 9521
rect 41931 9472 41932 9512
rect 41972 9472 41973 9512
rect 41931 9463 41973 9472
rect 42115 9512 42173 9513
rect 42115 9472 42124 9512
rect 42164 9472 42173 9512
rect 42115 9471 42173 9472
rect 42219 9512 42261 9521
rect 42219 9472 42220 9512
rect 42260 9472 42261 9512
rect 42219 9463 42261 9472
rect 42411 9512 42453 9521
rect 42411 9472 42412 9512
rect 42452 9472 42453 9512
rect 42411 9463 42453 9472
rect 42603 9512 42645 9521
rect 42603 9472 42604 9512
rect 42644 9472 42645 9512
rect 42603 9463 42645 9472
rect 42699 9512 42741 9521
rect 42699 9472 42700 9512
rect 42740 9472 42741 9512
rect 42699 9463 42741 9472
rect 42795 9512 42837 9521
rect 42795 9472 42796 9512
rect 42836 9472 42837 9512
rect 42795 9463 42837 9472
rect 42891 9512 42933 9521
rect 42891 9472 42892 9512
rect 42932 9472 42933 9512
rect 42891 9463 42933 9472
rect 45859 9512 45917 9513
rect 45859 9472 45868 9512
rect 45908 9472 45917 9512
rect 45859 9471 45917 9472
rect 46059 9512 46101 9521
rect 46059 9472 46060 9512
rect 46100 9472 46101 9512
rect 46059 9463 46101 9472
rect 46539 9512 46581 9521
rect 46539 9472 46540 9512
rect 46580 9472 46581 9512
rect 46539 9463 46581 9472
rect 46635 9512 46677 9521
rect 46635 9472 46636 9512
rect 46676 9472 46677 9512
rect 46635 9463 46677 9472
rect 46915 9512 46973 9513
rect 46915 9472 46924 9512
rect 46964 9472 46973 9512
rect 46915 9471 46973 9472
rect 50659 9512 50717 9513
rect 50659 9472 50668 9512
rect 50708 9472 50717 9512
rect 50659 9471 50717 9472
rect 52971 9512 53013 9521
rect 52971 9472 52972 9512
rect 53012 9472 53013 9512
rect 52971 9463 53013 9472
rect 53163 9512 53205 9521
rect 53163 9472 53164 9512
rect 53204 9472 53205 9512
rect 53731 9512 53789 9513
rect 53163 9463 53205 9472
rect 53261 9493 53319 9494
rect 53261 9453 53270 9493
rect 53310 9453 53319 9493
rect 53731 9472 53740 9512
rect 53780 9472 53789 9512
rect 53731 9471 53789 9472
rect 53931 9512 53973 9521
rect 53931 9472 53932 9512
rect 53972 9472 53973 9512
rect 53931 9463 53973 9472
rect 54219 9512 54261 9521
rect 54219 9472 54220 9512
rect 54260 9472 54261 9512
rect 54219 9463 54261 9472
rect 54403 9512 54461 9513
rect 54403 9472 54412 9512
rect 54452 9472 54461 9512
rect 54403 9471 54461 9472
rect 57771 9512 57813 9521
rect 57771 9472 57772 9512
rect 57812 9472 57813 9512
rect 57771 9463 57813 9472
rect 57963 9512 58005 9521
rect 57963 9472 57964 9512
rect 58004 9472 58005 9512
rect 57963 9463 58005 9472
rect 58051 9512 58109 9513
rect 58051 9472 58060 9512
rect 58100 9472 58109 9512
rect 58051 9471 58109 9472
rect 58339 9512 58397 9513
rect 58339 9472 58348 9512
rect 58388 9472 58397 9512
rect 58339 9471 58397 9472
rect 58635 9512 58677 9521
rect 58635 9472 58636 9512
rect 58676 9472 58677 9512
rect 58635 9463 58677 9472
rect 58731 9512 58773 9521
rect 58731 9472 58732 9512
rect 58772 9472 58773 9512
rect 58731 9463 58773 9472
rect 59595 9512 59637 9521
rect 59595 9472 59596 9512
rect 59636 9472 59637 9512
rect 59595 9463 59637 9472
rect 59971 9512 60029 9513
rect 59971 9472 59980 9512
rect 60020 9472 60029 9512
rect 59971 9471 60029 9472
rect 60835 9512 60893 9513
rect 60835 9472 60844 9512
rect 60884 9472 60893 9512
rect 60835 9471 60893 9472
rect 62563 9512 62621 9513
rect 62563 9472 62572 9512
rect 62612 9472 62621 9512
rect 62563 9471 62621 9472
rect 63427 9512 63485 9513
rect 63427 9472 63436 9512
rect 63476 9472 63485 9512
rect 63427 9471 63485 9472
rect 64779 9512 64821 9521
rect 64779 9472 64780 9512
rect 64820 9472 64821 9512
rect 64779 9463 64821 9472
rect 64971 9512 65013 9521
rect 64971 9472 64972 9512
rect 65012 9472 65013 9512
rect 64971 9463 65013 9472
rect 65059 9512 65117 9513
rect 65059 9472 65068 9512
rect 65108 9472 65117 9512
rect 65059 9471 65117 9472
rect 65251 9512 65309 9513
rect 65251 9472 65260 9512
rect 65300 9472 65309 9512
rect 65251 9471 65309 9472
rect 65451 9512 65493 9521
rect 65451 9472 65452 9512
rect 65492 9472 65493 9512
rect 65451 9463 65493 9472
rect 67267 9512 67325 9513
rect 67267 9472 67276 9512
rect 67316 9472 67325 9512
rect 67267 9471 67325 9472
rect 68131 9512 68189 9513
rect 68131 9472 68140 9512
rect 68180 9472 68189 9512
rect 68131 9471 68189 9472
rect 69867 9512 69909 9521
rect 69867 9472 69868 9512
rect 69908 9472 69909 9512
rect 69867 9463 69909 9472
rect 70059 9512 70101 9521
rect 70059 9472 70060 9512
rect 70100 9472 70101 9512
rect 70059 9463 70101 9472
rect 70147 9512 70205 9513
rect 70147 9472 70156 9512
rect 70196 9472 70205 9512
rect 70147 9471 70205 9472
rect 70723 9512 70781 9513
rect 70723 9472 70732 9512
rect 70772 9472 70781 9512
rect 70723 9471 70781 9472
rect 70827 9512 70869 9521
rect 70827 9472 70828 9512
rect 70868 9472 70869 9512
rect 70827 9463 70869 9472
rect 70923 9512 70965 9521
rect 70923 9472 70924 9512
rect 70964 9472 70965 9512
rect 70923 9463 70965 9472
rect 71299 9512 71357 9513
rect 71299 9472 71308 9512
rect 71348 9472 71357 9512
rect 71299 9471 71357 9472
rect 71499 9512 71541 9521
rect 71499 9472 71500 9512
rect 71540 9472 71541 9512
rect 71499 9463 71541 9472
rect 71683 9512 71741 9513
rect 71683 9472 71692 9512
rect 71732 9472 71741 9512
rect 71683 9471 71741 9472
rect 71883 9512 71925 9521
rect 71883 9472 71884 9512
rect 71924 9472 71925 9512
rect 71883 9463 71925 9472
rect 75627 9512 75669 9521
rect 75627 9472 75628 9512
rect 75668 9472 75669 9512
rect 75723 9493 75724 9533
rect 75764 9493 75765 9533
rect 75723 9484 75765 9493
rect 75819 9533 75861 9542
rect 75819 9493 75820 9533
rect 75860 9493 75861 9533
rect 76203 9525 76245 9534
rect 75819 9484 75861 9493
rect 76011 9512 76053 9521
rect 75627 9463 75669 9472
rect 76011 9472 76012 9512
rect 76052 9472 76053 9512
rect 76203 9485 76204 9525
rect 76244 9485 76245 9525
rect 76203 9476 76245 9485
rect 76291 9512 76349 9513
rect 76011 9463 76053 9472
rect 76291 9472 76300 9512
rect 76340 9472 76349 9512
rect 76291 9471 76349 9472
rect 77067 9512 77109 9521
rect 77067 9472 77068 9512
rect 77108 9472 77109 9512
rect 77067 9463 77109 9472
rect 77259 9512 77301 9521
rect 77259 9472 77260 9512
rect 77300 9472 77301 9512
rect 77259 9463 77301 9472
rect 77347 9512 77405 9513
rect 77347 9472 77356 9512
rect 77396 9472 77405 9512
rect 77347 9471 77405 9472
rect 77539 9512 77597 9513
rect 77539 9472 77548 9512
rect 77588 9472 77597 9512
rect 77539 9471 77597 9472
rect 77739 9512 77781 9521
rect 77739 9472 77740 9512
rect 77780 9472 77781 9512
rect 77739 9463 77781 9472
rect 77923 9512 77981 9513
rect 77923 9472 77932 9512
rect 77972 9472 77981 9512
rect 77923 9471 77981 9472
rect 78123 9512 78165 9521
rect 78123 9472 78124 9512
rect 78164 9472 78165 9512
rect 78123 9463 78165 9472
rect 53261 9452 53319 9453
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 1699 9428 1757 9429
rect 1699 9388 1708 9428
rect 1748 9388 1757 9428
rect 1699 9387 1757 9388
rect 52099 9428 52157 9429
rect 52099 9388 52108 9428
rect 52148 9388 52157 9428
rect 52099 9387 52157 9388
rect 57379 9428 57437 9429
rect 57379 9388 57388 9428
rect 57428 9388 57437 9428
rect 57379 9387 57437 9388
rect 59395 9428 59453 9429
rect 59395 9388 59404 9428
rect 59444 9388 59453 9428
rect 70339 9428 70397 9429
rect 59395 9387 59453 9388
rect 69465 9425 69523 9426
rect 3523 9386 3581 9387
rect 1323 9344 1365 9353
rect 3523 9346 3532 9386
rect 3572 9346 3581 9386
rect 69465 9385 69474 9425
rect 69514 9385 69523 9425
rect 70339 9388 70348 9428
rect 70388 9388 70397 9428
rect 70339 9387 70397 9388
rect 76483 9428 76541 9429
rect 76483 9388 76492 9428
rect 76532 9388 76541 9428
rect 76483 9387 76541 9388
rect 69465 9384 69523 9385
rect 3523 9345 3581 9346
rect 1323 9304 1324 9344
rect 1364 9304 1365 9344
rect 1323 9295 1365 9304
rect 39435 9344 39477 9353
rect 39435 9304 39436 9344
rect 39476 9304 39477 9344
rect 39435 9295 39477 9304
rect 41451 9344 41493 9353
rect 41451 9304 41452 9344
rect 41492 9304 41493 9344
rect 41451 9295 41493 9304
rect 41931 9344 41973 9353
rect 41931 9304 41932 9344
rect 41972 9304 41973 9344
rect 41931 9295 41973 9304
rect 44715 9344 44757 9353
rect 44715 9304 44716 9344
rect 44756 9304 44757 9344
rect 44715 9295 44757 9304
rect 46243 9344 46301 9345
rect 46243 9304 46252 9344
rect 46292 9304 46301 9344
rect 46243 9303 46301 9304
rect 47211 9344 47253 9353
rect 47211 9304 47212 9344
rect 47252 9304 47253 9344
rect 47211 9295 47253 9304
rect 50379 9344 50421 9353
rect 50379 9304 50380 9344
rect 50420 9304 50421 9344
rect 50379 9295 50421 9304
rect 54891 9344 54933 9353
rect 54891 9304 54892 9344
rect 54932 9304 54933 9344
rect 54891 9295 54933 9304
rect 56427 9344 56469 9353
rect 56427 9304 56428 9344
rect 56468 9304 56469 9344
rect 56427 9295 56469 9304
rect 69867 9344 69909 9353
rect 69867 9304 69868 9344
rect 69908 9304 69909 9344
rect 69867 9295 69909 9304
rect 72171 9344 72213 9353
rect 72171 9304 72172 9344
rect 72212 9304 72213 9344
rect 72171 9295 72213 9304
rect 73899 9344 73941 9353
rect 73899 9304 73900 9344
rect 73940 9304 73941 9344
rect 73899 9295 73941 9304
rect 76011 9344 76053 9353
rect 76011 9304 76012 9344
rect 76052 9304 76053 9344
rect 76011 9295 76053 9304
rect 77643 9344 77685 9353
rect 77643 9304 77644 9344
rect 77684 9304 77685 9344
rect 77643 9295 77685 9304
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 3819 9260 3861 9269
rect 3819 9220 3820 9260
rect 3860 9220 3861 9260
rect 3819 9211 3861 9220
rect 7171 9260 7229 9261
rect 7171 9220 7180 9260
rect 7220 9220 7229 9260
rect 7171 9219 7229 9220
rect 42411 9260 42453 9269
rect 42411 9220 42412 9260
rect 42452 9220 42453 9260
rect 42411 9211 42453 9220
rect 45963 9260 46005 9269
rect 45963 9220 45964 9260
rect 46004 9220 46005 9260
rect 45963 9211 46005 9220
rect 52683 9260 52725 9269
rect 52683 9220 52684 9260
rect 52724 9220 52725 9260
rect 52683 9211 52725 9220
rect 53835 9260 53877 9269
rect 53835 9220 53836 9260
rect 53876 9220 53877 9260
rect 53835 9211 53877 9220
rect 54315 9260 54357 9269
rect 54315 9220 54316 9260
rect 54356 9220 54357 9260
rect 54315 9211 54357 9220
rect 57579 9260 57621 9269
rect 57579 9220 57580 9260
rect 57620 9220 57621 9260
rect 57579 9211 57621 9220
rect 57771 9260 57813 9269
rect 57771 9220 57772 9260
rect 57812 9220 57813 9260
rect 57771 9211 57813 9220
rect 59011 9260 59069 9261
rect 59011 9220 59020 9260
rect 59060 9220 59069 9260
rect 59011 9219 59069 9220
rect 59211 9260 59253 9269
rect 59211 9220 59212 9260
rect 59252 9220 59253 9260
rect 59211 9211 59253 9220
rect 61987 9260 62045 9261
rect 61987 9220 61996 9260
rect 62036 9220 62045 9260
rect 61987 9219 62045 9220
rect 64579 9260 64637 9261
rect 64579 9220 64588 9260
rect 64628 9220 64637 9260
rect 64579 9219 64637 9220
rect 69283 9260 69341 9261
rect 69283 9220 69292 9260
rect 69332 9220 69341 9260
rect 69283 9219 69341 9220
rect 69675 9260 69717 9269
rect 69675 9220 69676 9260
rect 69716 9220 69717 9260
rect 69675 9211 69717 9220
rect 70539 9260 70581 9269
rect 70539 9220 70540 9260
rect 70580 9220 70581 9260
rect 70539 9211 70581 9220
rect 71403 9260 71445 9269
rect 71403 9220 71404 9260
rect 71444 9220 71445 9260
rect 71403 9211 71445 9220
rect 71787 9260 71829 9269
rect 71787 9220 71788 9260
rect 71828 9220 71829 9260
rect 71787 9211 71829 9220
rect 76683 9260 76725 9269
rect 76683 9220 76684 9260
rect 76724 9220 76725 9260
rect 76683 9211 76725 9220
rect 78027 9260 78069 9269
rect 78027 9220 78028 9260
rect 78068 9220 78069 9260
rect 78027 9211 78069 9220
rect 576 9092 79584 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 75112 9092
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75480 9052 79584 9092
rect 576 9028 79584 9052
rect 43939 8924 43997 8925
rect 43939 8884 43948 8924
rect 43988 8884 43997 8924
rect 43939 8883 43997 8884
rect 46627 8924 46685 8925
rect 46627 8884 46636 8924
rect 46676 8884 46685 8924
rect 46627 8883 46685 8884
rect 51339 8924 51381 8933
rect 51339 8884 51340 8924
rect 51380 8884 51381 8924
rect 51339 8875 51381 8884
rect 53923 8924 53981 8925
rect 53923 8884 53932 8924
rect 53972 8884 53981 8924
rect 53923 8883 53981 8884
rect 56803 8924 56861 8925
rect 56803 8884 56812 8924
rect 56852 8884 56861 8924
rect 56803 8883 56861 8884
rect 69771 8924 69813 8933
rect 69771 8884 69772 8924
rect 69812 8884 69813 8924
rect 69771 8875 69813 8884
rect 71491 8924 71549 8925
rect 71491 8884 71500 8924
rect 71540 8884 71549 8924
rect 71491 8883 71549 8884
rect 74083 8924 74141 8925
rect 74083 8884 74092 8924
rect 74132 8884 74141 8924
rect 74083 8883 74141 8884
rect 79459 8924 79517 8925
rect 79459 8884 79468 8924
rect 79508 8884 79517 8924
rect 79459 8883 79517 8884
rect 49323 8840 49365 8849
rect 49323 8800 49324 8840
rect 49364 8800 49365 8840
rect 58923 8840 58965 8849
rect 49323 8791 49365 8800
rect 50955 8798 50997 8807
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 3531 8756 3573 8765
rect 3531 8716 3532 8756
rect 3572 8716 3573 8756
rect 50955 8758 50956 8798
rect 50996 8758 50997 8798
rect 58923 8800 58924 8840
rect 58964 8800 58965 8840
rect 58923 8791 58965 8800
rect 60939 8840 60981 8849
rect 60939 8800 60940 8840
rect 60980 8800 60981 8840
rect 60939 8791 60981 8800
rect 66507 8840 66549 8849
rect 66507 8800 66508 8840
rect 66548 8800 66549 8840
rect 66507 8791 66549 8800
rect 68523 8840 68565 8849
rect 68523 8800 68524 8840
rect 68564 8800 68565 8840
rect 68523 8791 68565 8800
rect 69195 8840 69237 8849
rect 69195 8800 69196 8840
rect 69236 8800 69237 8840
rect 69195 8791 69237 8800
rect 70059 8840 70101 8849
rect 70059 8800 70060 8840
rect 70100 8800 70101 8840
rect 70059 8791 70101 8800
rect 74283 8840 74325 8849
rect 74283 8800 74284 8840
rect 74324 8800 74325 8840
rect 74283 8791 74325 8800
rect 76867 8840 76925 8841
rect 76867 8800 76876 8840
rect 76916 8800 76925 8840
rect 76867 8799 76925 8800
rect 50955 8749 50997 8758
rect 58243 8756 58301 8757
rect 3531 8707 3573 8716
rect 58243 8716 58252 8756
rect 58292 8716 58301 8756
rect 58243 8715 58301 8716
rect 58723 8756 58781 8757
rect 58723 8716 58732 8756
rect 58772 8716 58781 8756
rect 58723 8715 58781 8716
rect 59691 8756 59733 8765
rect 59691 8716 59692 8756
rect 59732 8716 59733 8756
rect 59691 8707 59733 8716
rect 64771 8756 64829 8757
rect 64771 8716 64780 8756
rect 64820 8716 64829 8756
rect 64771 8715 64829 8716
rect 70243 8756 70301 8757
rect 70243 8716 70252 8756
rect 70292 8716 70301 8756
rect 70243 8715 70301 8716
rect 53251 8689 53309 8690
rect 1507 8672 1565 8673
rect 1507 8632 1516 8672
rect 1556 8632 1565 8672
rect 1507 8631 1565 8632
rect 2371 8672 2429 8673
rect 2371 8632 2380 8672
rect 2420 8632 2429 8672
rect 2371 8631 2429 8632
rect 4771 8672 4829 8673
rect 4771 8632 4780 8672
rect 4820 8632 4829 8672
rect 4771 8631 4829 8632
rect 4971 8672 5013 8681
rect 4971 8632 4972 8672
rect 5012 8632 5013 8672
rect 4971 8623 5013 8632
rect 41923 8672 41981 8673
rect 41923 8632 41932 8672
rect 41972 8632 41981 8672
rect 41923 8631 41981 8632
rect 42787 8672 42845 8673
rect 42787 8632 42796 8672
rect 42836 8632 42845 8672
rect 42787 8631 42845 8632
rect 44611 8672 44669 8673
rect 44611 8632 44620 8672
rect 44660 8632 44669 8672
rect 44611 8631 44669 8632
rect 45475 8672 45533 8673
rect 45475 8632 45484 8672
rect 45524 8632 45533 8672
rect 45475 8631 45533 8632
rect 48451 8672 48509 8673
rect 48451 8632 48460 8672
rect 48500 8632 48509 8672
rect 48451 8631 48509 8632
rect 48651 8672 48693 8681
rect 48651 8632 48652 8672
rect 48692 8632 48693 8672
rect 48651 8623 48693 8632
rect 48843 8672 48885 8681
rect 48843 8632 48844 8672
rect 48884 8632 48885 8672
rect 48843 8623 48885 8632
rect 49035 8672 49077 8681
rect 49035 8632 49036 8672
rect 49076 8632 49077 8672
rect 49035 8623 49077 8632
rect 49123 8672 49181 8673
rect 49123 8632 49132 8672
rect 49172 8632 49181 8672
rect 49123 8631 49181 8632
rect 49699 8672 49757 8673
rect 49699 8632 49708 8672
rect 49748 8632 49757 8672
rect 49699 8631 49757 8632
rect 49803 8672 49845 8681
rect 49803 8632 49804 8672
rect 49844 8632 49845 8672
rect 49803 8623 49845 8632
rect 49899 8672 49941 8681
rect 49899 8632 49900 8672
rect 49940 8632 49941 8672
rect 49899 8623 49941 8632
rect 51339 8672 51381 8681
rect 51339 8632 51340 8672
rect 51380 8632 51381 8672
rect 51339 8623 51381 8632
rect 51531 8672 51573 8681
rect 51531 8632 51532 8672
rect 51572 8632 51573 8672
rect 51531 8623 51573 8632
rect 51619 8672 51677 8673
rect 51619 8632 51628 8672
rect 51668 8632 51677 8672
rect 51619 8631 51677 8632
rect 52203 8672 52245 8681
rect 52203 8632 52204 8672
rect 52244 8632 52245 8672
rect 52203 8623 52245 8632
rect 52299 8672 52341 8681
rect 52299 8632 52300 8672
rect 52340 8632 52341 8672
rect 52299 8623 52341 8632
rect 52395 8672 52437 8681
rect 52395 8632 52396 8672
rect 52436 8632 52437 8672
rect 52395 8623 52437 8632
rect 52491 8672 52533 8681
rect 52491 8632 52492 8672
rect 52532 8632 52533 8672
rect 52491 8623 52533 8632
rect 52683 8672 52725 8681
rect 52683 8632 52684 8672
rect 52724 8632 52725 8672
rect 52683 8623 52725 8632
rect 52875 8672 52917 8681
rect 52875 8632 52876 8672
rect 52916 8632 52917 8672
rect 52875 8623 52917 8632
rect 52963 8672 53021 8673
rect 52963 8632 52972 8672
rect 53012 8632 53021 8672
rect 53251 8649 53260 8689
rect 53300 8649 53309 8689
rect 53251 8648 53309 8649
rect 53547 8672 53589 8681
rect 52963 8631 53021 8632
rect 53547 8632 53548 8672
rect 53588 8632 53589 8672
rect 53547 8623 53589 8632
rect 54787 8672 54845 8673
rect 54787 8632 54796 8672
rect 54836 8632 54845 8672
rect 54787 8631 54845 8632
rect 55651 8672 55709 8673
rect 55651 8632 55660 8672
rect 55700 8632 55709 8672
rect 55651 8631 55709 8632
rect 57771 8672 57813 8681
rect 57771 8632 57772 8672
rect 57812 8632 57813 8672
rect 57771 8623 57813 8632
rect 57867 8672 57909 8681
rect 57867 8632 57868 8672
rect 57908 8632 57909 8672
rect 57867 8623 57909 8632
rect 57963 8672 58005 8681
rect 57963 8632 57964 8672
rect 58004 8632 58005 8672
rect 57963 8623 58005 8632
rect 58059 8672 58101 8681
rect 58059 8632 58060 8672
rect 58100 8632 58101 8672
rect 58059 8623 58101 8632
rect 59115 8672 59157 8681
rect 59115 8632 59116 8672
rect 59156 8632 59157 8672
rect 59115 8623 59157 8632
rect 59307 8672 59349 8681
rect 59307 8632 59308 8672
rect 59348 8632 59349 8672
rect 59307 8623 59349 8632
rect 59395 8672 59453 8673
rect 59395 8632 59404 8672
rect 59444 8632 59453 8672
rect 59395 8631 59453 8632
rect 59595 8672 59637 8681
rect 59595 8632 59596 8672
rect 59636 8632 59637 8672
rect 59595 8623 59637 8632
rect 59779 8672 59837 8673
rect 59779 8632 59788 8672
rect 59828 8632 59837 8672
rect 59779 8631 59837 8632
rect 59971 8672 60029 8673
rect 59971 8632 59980 8672
rect 60020 8632 60029 8672
rect 59971 8631 60029 8632
rect 60075 8672 60117 8681
rect 60075 8632 60076 8672
rect 60116 8632 60117 8672
rect 60075 8623 60117 8632
rect 60171 8672 60213 8681
rect 60171 8632 60172 8672
rect 60212 8632 60213 8672
rect 60171 8623 60213 8632
rect 63819 8672 63861 8681
rect 63819 8632 63820 8672
rect 63860 8632 63861 8672
rect 63819 8623 63861 8632
rect 63915 8672 63957 8681
rect 63915 8632 63916 8672
rect 63956 8632 63957 8672
rect 63915 8623 63957 8632
rect 64011 8672 64053 8681
rect 64011 8632 64012 8672
rect 64052 8632 64053 8672
rect 64011 8623 64053 8632
rect 64107 8672 64149 8681
rect 64107 8632 64108 8672
rect 64148 8632 64149 8672
rect 64107 8623 64149 8632
rect 64299 8672 64341 8681
rect 64299 8632 64300 8672
rect 64340 8632 64341 8672
rect 64299 8623 64341 8632
rect 64491 8672 64533 8681
rect 64491 8632 64492 8672
rect 64532 8632 64533 8672
rect 64491 8623 64533 8632
rect 64579 8672 64637 8673
rect 64579 8632 64588 8672
rect 64628 8632 64637 8672
rect 64579 8631 64637 8632
rect 68715 8672 68757 8681
rect 68715 8632 68716 8672
rect 68756 8632 68757 8672
rect 68715 8623 68757 8632
rect 68907 8672 68949 8681
rect 68907 8632 68908 8672
rect 68948 8632 68949 8672
rect 68907 8623 68949 8632
rect 68995 8672 69053 8673
rect 68995 8632 69004 8672
rect 69044 8632 69053 8672
rect 68995 8631 69053 8632
rect 69195 8672 69237 8681
rect 69195 8632 69196 8672
rect 69236 8632 69237 8672
rect 69195 8623 69237 8632
rect 69387 8672 69429 8681
rect 69387 8632 69388 8672
rect 69428 8632 69429 8672
rect 69387 8623 69429 8632
rect 69475 8672 69533 8673
rect 69475 8632 69484 8672
rect 69524 8632 69533 8672
rect 69867 8672 69909 8681
rect 69475 8631 69533 8632
rect 69667 8651 69725 8652
rect 69667 8611 69676 8651
rect 69716 8611 69725 8651
rect 69867 8632 69868 8672
rect 69908 8632 69909 8672
rect 69867 8623 69909 8632
rect 70819 8672 70877 8673
rect 70819 8632 70828 8672
rect 70868 8632 70877 8672
rect 70819 8631 70877 8632
rect 71115 8672 71157 8681
rect 71115 8632 71116 8672
rect 71156 8632 71157 8672
rect 71115 8623 71157 8632
rect 72067 8672 72125 8673
rect 72067 8632 72076 8672
rect 72116 8632 72125 8672
rect 72067 8631 72125 8632
rect 72931 8672 72989 8673
rect 72931 8632 72940 8672
rect 72980 8632 72989 8672
rect 72931 8631 72989 8632
rect 75627 8672 75669 8681
rect 75627 8632 75628 8672
rect 75668 8632 75669 8672
rect 75627 8623 75669 8632
rect 75819 8672 75861 8681
rect 75819 8632 75820 8672
rect 75860 8632 75861 8672
rect 75819 8623 75861 8632
rect 75907 8672 75965 8673
rect 75907 8632 75916 8672
rect 75956 8632 75965 8672
rect 75907 8631 75965 8632
rect 76195 8672 76253 8673
rect 76195 8632 76204 8672
rect 76244 8632 76253 8672
rect 76195 8631 76253 8632
rect 76491 8672 76533 8681
rect 76491 8632 76492 8672
rect 76532 8632 76533 8672
rect 76491 8623 76533 8632
rect 77443 8672 77501 8673
rect 77443 8632 77452 8672
rect 77492 8632 77501 8672
rect 77443 8631 77501 8632
rect 78307 8672 78365 8673
rect 78307 8632 78316 8672
rect 78356 8632 78365 8672
rect 78307 8631 78365 8632
rect 69667 8610 69725 8611
rect 1131 8588 1173 8597
rect 1131 8548 1132 8588
rect 1172 8548 1173 8588
rect 1131 8539 1173 8548
rect 4875 8588 4917 8597
rect 4875 8548 4876 8588
rect 4916 8548 4917 8588
rect 4875 8539 4917 8548
rect 41547 8588 41589 8597
rect 41547 8548 41548 8588
rect 41588 8548 41589 8588
rect 41547 8539 41589 8548
rect 44235 8588 44277 8597
rect 44235 8548 44236 8588
rect 44276 8548 44277 8588
rect 44235 8539 44277 8548
rect 48555 8588 48597 8597
rect 48555 8548 48556 8588
rect 48596 8548 48597 8588
rect 48555 8539 48597 8548
rect 53643 8588 53685 8597
rect 53643 8548 53644 8588
rect 53684 8548 53685 8588
rect 53643 8539 53685 8548
rect 54411 8588 54453 8597
rect 54411 8548 54412 8588
rect 54452 8548 54453 8588
rect 54411 8539 54453 8548
rect 59211 8588 59253 8597
rect 59211 8548 59212 8588
rect 59252 8548 59253 8588
rect 59211 8539 59253 8548
rect 64395 8588 64437 8597
rect 64395 8548 64396 8588
rect 64436 8548 64437 8588
rect 64395 8539 64437 8548
rect 71211 8588 71253 8597
rect 71211 8548 71212 8588
rect 71252 8548 71253 8588
rect 71211 8539 71253 8548
rect 71691 8588 71733 8597
rect 71691 8548 71692 8588
rect 71732 8548 71733 8588
rect 71691 8539 71733 8548
rect 75723 8588 75765 8597
rect 75723 8548 75724 8588
rect 75764 8548 75765 8588
rect 75723 8539 75765 8548
rect 76587 8588 76629 8597
rect 76587 8548 76588 8588
rect 76628 8548 76629 8588
rect 76587 8539 76629 8548
rect 77067 8588 77109 8597
rect 77067 8548 77068 8588
rect 77108 8548 77109 8588
rect 77067 8539 77109 8548
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 43939 8504 43997 8505
rect 43939 8464 43948 8504
rect 43988 8464 43997 8504
rect 43939 8463 43997 8464
rect 46627 8504 46685 8505
rect 46627 8464 46636 8504
rect 46676 8464 46685 8504
rect 46627 8463 46685 8464
rect 48931 8504 48989 8505
rect 48931 8464 48940 8504
rect 48980 8464 48989 8504
rect 48931 8463 48989 8464
rect 52771 8504 52829 8505
rect 52771 8464 52780 8504
rect 52820 8464 52829 8504
rect 52771 8463 52829 8464
rect 58443 8504 58485 8513
rect 58443 8464 58444 8504
rect 58484 8464 58485 8504
rect 58443 8455 58485 8464
rect 64971 8504 65013 8513
rect 64971 8464 64972 8504
rect 65012 8464 65013 8504
rect 64971 8455 65013 8464
rect 68803 8504 68861 8505
rect 68803 8464 68812 8504
rect 68852 8464 68861 8504
rect 68803 8463 68861 8464
rect 576 8336 79584 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 76352 8336
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76720 8296 79584 8336
rect 576 8272 79584 8296
rect 2371 8168 2429 8169
rect 2371 8128 2380 8168
rect 2420 8128 2429 8168
rect 2371 8127 2429 8128
rect 4675 8168 4733 8169
rect 4675 8128 4684 8168
rect 4724 8128 4733 8168
rect 4675 8127 4733 8128
rect 7459 8168 7517 8169
rect 7459 8128 7468 8168
rect 7508 8128 7517 8168
rect 7459 8127 7517 8128
rect 44995 8168 45053 8169
rect 44995 8128 45004 8168
rect 45044 8128 45053 8168
rect 44995 8127 45053 8128
rect 52867 8168 52925 8169
rect 52867 8128 52876 8168
rect 52916 8128 52925 8168
rect 52867 8127 52925 8128
rect 58339 8168 58397 8169
rect 58339 8128 58348 8168
rect 58388 8128 58397 8168
rect 58339 8127 58397 8128
rect 62851 8168 62909 8169
rect 62851 8128 62860 8168
rect 62900 8128 62909 8168
rect 62851 8127 62909 8128
rect 64099 8168 64157 8169
rect 64099 8128 64108 8168
rect 64148 8128 64157 8168
rect 64099 8127 64157 8128
rect 65635 8168 65693 8169
rect 65635 8128 65644 8168
rect 65684 8128 65693 8168
rect 65635 8127 65693 8128
rect 68419 8168 68477 8169
rect 68419 8128 68428 8168
rect 68468 8128 68477 8168
rect 68419 8127 68477 8128
rect 71011 8168 71069 8169
rect 71011 8128 71020 8168
rect 71060 8128 71069 8168
rect 71011 8127 71069 8128
rect 71491 8168 71549 8169
rect 71491 8128 71500 8168
rect 71540 8128 71549 8168
rect 71491 8127 71549 8128
rect 75907 8168 75965 8169
rect 75907 8128 75916 8168
rect 75956 8128 75965 8168
rect 75907 8127 75965 8128
rect 77059 8168 77117 8169
rect 77059 8128 77068 8168
rect 77108 8128 77117 8168
rect 77059 8127 77117 8128
rect 5067 8084 5109 8093
rect 5067 8044 5068 8084
rect 5108 8044 5109 8084
rect 5067 8035 5109 8044
rect 54123 8084 54165 8093
rect 54123 8044 54124 8084
rect 54164 8044 54165 8084
rect 54123 8035 54165 8044
rect 55947 8084 55989 8093
rect 55947 8044 55948 8084
rect 55988 8044 55989 8084
rect 55947 8035 55989 8044
rect 66027 8084 66069 8093
rect 66027 8044 66028 8084
rect 66068 8044 66069 8084
rect 66027 8035 66069 8044
rect 68619 8084 68661 8093
rect 68619 8044 68620 8084
rect 68660 8044 68661 8084
rect 68619 8035 68661 8044
rect 53259 8021 53301 8030
rect 1803 8000 1845 8009
rect 1803 7960 1804 8000
rect 1844 7960 1845 8000
rect 1803 7951 1845 7960
rect 1899 8000 1941 8009
rect 1899 7960 1900 8000
rect 1940 7960 1941 8000
rect 1899 7951 1941 7960
rect 1995 8000 2037 8009
rect 1995 7960 1996 8000
rect 2036 7960 2037 8000
rect 1995 7951 2037 7960
rect 2091 8000 2133 8009
rect 2091 7960 2092 8000
rect 2132 7960 2133 8000
rect 2091 7951 2133 7960
rect 2283 8000 2325 8009
rect 2283 7960 2284 8000
rect 2324 7960 2325 8000
rect 2283 7951 2325 7960
rect 2475 8000 2517 8009
rect 2475 7960 2476 8000
rect 2516 7960 2517 8000
rect 2475 7951 2517 7960
rect 2563 8000 2621 8001
rect 2563 7960 2572 8000
rect 2612 7960 2621 8000
rect 2563 7959 2621 7960
rect 2763 8000 2805 8009
rect 2763 7960 2764 8000
rect 2804 7960 2805 8000
rect 2763 7951 2805 7960
rect 2955 8000 2997 8009
rect 2955 7960 2956 8000
rect 2996 7960 2997 8000
rect 2955 7951 2997 7960
rect 3043 8000 3101 8001
rect 3043 7960 3052 8000
rect 3092 7960 3101 8000
rect 3043 7959 3101 7960
rect 3427 8000 3485 8001
rect 3427 7960 3436 8000
rect 3476 7960 3485 8000
rect 3427 7959 3485 7960
rect 3723 8000 3765 8009
rect 3723 7960 3724 8000
rect 3764 7960 3765 8000
rect 3723 7951 3765 7960
rect 3819 8000 3861 8009
rect 3819 7960 3820 8000
rect 3860 7960 3861 8000
rect 3819 7951 3861 7960
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4779 8000 4821 8009
rect 4779 7960 4780 8000
rect 4820 7960 4821 8000
rect 4779 7951 4821 7960
rect 4867 8000 4925 8001
rect 4867 7960 4876 8000
rect 4916 7960 4925 8000
rect 4867 7959 4925 7960
rect 5443 8000 5501 8001
rect 5443 7960 5452 8000
rect 5492 7960 5501 8000
rect 5443 7959 5501 7960
rect 6307 8000 6365 8001
rect 6307 7960 6316 8000
rect 6356 7960 6365 8000
rect 6307 7959 6365 7960
rect 44131 8000 44189 8001
rect 44131 7960 44140 8000
rect 44180 7960 44189 8000
rect 44131 7959 44189 7960
rect 44235 8000 44277 8009
rect 44235 7960 44236 8000
rect 44276 7960 44277 8000
rect 44235 7951 44277 7960
rect 44427 8000 44469 8009
rect 44427 7960 44428 8000
rect 44468 7960 44469 8000
rect 44427 7951 44469 7960
rect 44803 8000 44861 8001
rect 44803 7960 44812 8000
rect 44852 7960 44861 8000
rect 44803 7959 44861 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 45099 8000 45141 8009
rect 45099 7960 45100 8000
rect 45140 7960 45141 8000
rect 45099 7951 45141 7960
rect 45387 8000 45429 8009
rect 45387 7960 45388 8000
rect 45428 7960 45429 8000
rect 45387 7951 45429 7960
rect 45483 8000 45525 8009
rect 45483 7960 45484 8000
rect 45524 7960 45525 8000
rect 45483 7951 45525 7960
rect 45579 8000 45621 8009
rect 45579 7960 45580 8000
rect 45620 7960 45621 8000
rect 45579 7951 45621 7960
rect 45675 8000 45717 8009
rect 45675 7960 45676 8000
rect 45716 7960 45717 8000
rect 45675 7951 45717 7960
rect 46723 8000 46781 8001
rect 46723 7960 46732 8000
rect 46772 7960 46781 8000
rect 46723 7959 46781 7960
rect 46827 8000 46869 8009
rect 46827 7960 46828 8000
rect 46868 7960 46869 8000
rect 46827 7951 46869 7960
rect 47019 8000 47061 8009
rect 47019 7960 47020 8000
rect 47060 7960 47061 8000
rect 47019 7951 47061 7960
rect 47203 8000 47261 8001
rect 47203 7960 47212 8000
rect 47252 7960 47261 8000
rect 47203 7959 47261 7960
rect 47307 8000 47349 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 47499 8000 47541 8009
rect 47499 7960 47500 8000
rect 47540 7960 47541 8000
rect 47499 7951 47541 7960
rect 47971 8000 48029 8001
rect 47971 7960 47980 8000
rect 48020 7960 48029 8000
rect 47971 7959 48029 7960
rect 48267 8000 48309 8009
rect 48267 7960 48268 8000
rect 48308 7960 48309 8000
rect 48267 7951 48309 7960
rect 48363 8000 48405 8009
rect 49219 8000 49277 8001
rect 48363 7960 48364 8000
rect 48404 7960 48405 8000
rect 48363 7951 48405 7960
rect 48835 7999 48893 8000
rect 48835 7959 48844 7999
rect 48884 7959 48893 7999
rect 49219 7960 49228 8000
rect 49268 7960 49277 8000
rect 49219 7959 49277 7960
rect 50179 8000 50237 8001
rect 50179 7960 50188 8000
rect 50228 7960 50237 8000
rect 50179 7959 50237 7960
rect 50475 8000 50517 8009
rect 50475 7960 50476 8000
rect 50516 7960 50517 8000
rect 48835 7958 48893 7959
rect 50475 7951 50517 7960
rect 50851 8000 50909 8001
rect 50851 7960 50860 8000
rect 50900 7960 50909 8000
rect 50851 7959 50909 7960
rect 51715 8000 51773 8001
rect 51715 7960 51724 8000
rect 51764 7960 51773 8000
rect 51715 7959 51773 7960
rect 53067 8000 53109 8009
rect 53067 7960 53068 8000
rect 53108 7960 53109 8000
rect 53067 7951 53109 7960
rect 53163 8000 53205 8009
rect 53163 7960 53164 8000
rect 53204 7960 53205 8000
rect 53259 7981 53260 8021
rect 53300 7981 53301 8021
rect 53259 7972 53301 7981
rect 53355 8000 53397 8009
rect 53163 7951 53205 7960
rect 53355 7960 53356 8000
rect 53396 7960 53397 8000
rect 53355 7951 53397 7960
rect 54027 8000 54069 8009
rect 54027 7960 54028 8000
rect 54068 7960 54069 8000
rect 54027 7951 54069 7960
rect 54219 8000 54261 8009
rect 54219 7960 54220 8000
rect 54260 7960 54261 8000
rect 54219 7951 54261 7960
rect 54307 8000 54365 8001
rect 54307 7960 54316 8000
rect 54356 7960 54365 8000
rect 54307 7959 54365 7960
rect 56323 8000 56381 8001
rect 56323 7960 56332 8000
rect 56372 7960 56381 8000
rect 56323 7959 56381 7960
rect 57187 8000 57245 8001
rect 57187 7960 57196 8000
rect 57236 7960 57245 8000
rect 57187 7959 57245 7960
rect 58531 8000 58589 8001
rect 58531 7960 58540 8000
rect 58580 7960 58589 8000
rect 58531 7959 58589 7960
rect 58635 8000 58677 8009
rect 58635 7960 58636 8000
rect 58676 7960 58677 8000
rect 58635 7951 58677 7960
rect 58827 8000 58869 8009
rect 58827 7960 58828 8000
rect 58868 7960 58869 8000
rect 58827 7951 58869 7960
rect 60075 8000 60117 8009
rect 60075 7960 60076 8000
rect 60116 7960 60117 8000
rect 60075 7951 60117 7960
rect 60259 8000 60317 8001
rect 60259 7960 60268 8000
rect 60308 7960 60317 8000
rect 60259 7959 60317 7960
rect 60459 8000 60501 8009
rect 60459 7960 60460 8000
rect 60500 7960 60501 8000
rect 60459 7951 60501 7960
rect 60835 8000 60893 8001
rect 60835 7960 60844 8000
rect 60884 7960 60893 8000
rect 60835 7959 60893 7960
rect 61699 8000 61757 8001
rect 61699 7960 61708 8000
rect 61748 7960 61757 8000
rect 61699 7959 61757 7960
rect 63627 8000 63669 8009
rect 63627 7960 63628 8000
rect 63668 7960 63669 8000
rect 63627 7951 63669 7960
rect 63819 8000 63861 8009
rect 63819 7960 63820 8000
rect 63860 7960 63861 8000
rect 63819 7951 63861 7960
rect 63907 8000 63965 8001
rect 63907 7960 63916 8000
rect 63956 7960 63965 8000
rect 63907 7959 63965 7960
rect 64203 8000 64245 8009
rect 64203 7960 64204 8000
rect 64244 7960 64245 8000
rect 64203 7951 64245 7960
rect 64299 8000 64341 8009
rect 64299 7960 64300 8000
rect 64340 7960 64341 8000
rect 64299 7951 64341 7960
rect 64395 8000 64437 8009
rect 64395 7960 64396 8000
rect 64436 7960 64437 8000
rect 64395 7951 64437 7960
rect 64675 8000 64733 8001
rect 64675 7960 64684 8000
rect 64724 7960 64733 8000
rect 64675 7959 64733 7960
rect 64971 8000 65013 8009
rect 64971 7960 64972 8000
rect 65012 7960 65013 8000
rect 64971 7951 65013 7960
rect 65067 8000 65109 8009
rect 65067 7960 65068 8000
rect 65108 7960 65109 8000
rect 65067 7951 65109 7960
rect 65547 8000 65589 8009
rect 65547 7960 65548 8000
rect 65588 7960 65589 8000
rect 65547 7951 65589 7960
rect 65739 8000 65781 8009
rect 65739 7960 65740 8000
rect 65780 7960 65781 8000
rect 65739 7951 65781 7960
rect 65827 8000 65885 8001
rect 65827 7960 65836 8000
rect 65876 7960 65885 8000
rect 65827 7959 65885 7960
rect 66403 8000 66461 8001
rect 66403 7960 66412 8000
rect 66452 7960 66461 8000
rect 66403 7959 66461 7960
rect 67267 8000 67325 8001
rect 67267 7960 67276 8000
rect 67316 7960 67325 8000
rect 67267 7959 67325 7960
rect 68995 8000 69053 8001
rect 68995 7960 69004 8000
rect 69044 7960 69053 8000
rect 68995 7959 69053 7960
rect 69859 8000 69917 8001
rect 69859 7960 69868 8000
rect 69908 7960 69917 8000
rect 69859 7959 69917 7960
rect 71403 8000 71445 8009
rect 71403 7960 71404 8000
rect 71444 7960 71445 8000
rect 71403 7951 71445 7960
rect 71595 8000 71637 8009
rect 71595 7960 71596 8000
rect 71636 7960 71637 8000
rect 71595 7951 71637 7960
rect 71683 8000 71741 8001
rect 71683 7960 71692 8000
rect 71732 7960 71741 8000
rect 71683 7959 71741 7960
rect 73515 8000 73557 8009
rect 73515 7960 73516 8000
rect 73556 7960 73557 8000
rect 73515 7951 73557 7960
rect 73891 8000 73949 8001
rect 73891 7960 73900 8000
rect 73940 7960 73949 8000
rect 73891 7959 73949 7960
rect 74755 8000 74813 8001
rect 74755 7960 74764 8000
rect 74804 7960 74813 8000
rect 74755 7959 74813 7960
rect 76107 8000 76149 8009
rect 76107 7960 76108 8000
rect 76148 7960 76149 8000
rect 76107 7951 76149 7960
rect 76203 8000 76245 8009
rect 76203 7960 76204 8000
rect 76244 7960 76245 8000
rect 76203 7951 76245 7960
rect 76299 8000 76341 8009
rect 76299 7960 76300 8000
rect 76340 7960 76341 8000
rect 76299 7951 76341 7960
rect 76395 8000 76437 8009
rect 76395 7960 76396 8000
rect 76436 7960 76437 8000
rect 76395 7951 76437 7960
rect 76579 8000 76637 8001
rect 76579 7960 76588 8000
rect 76628 7960 76637 8000
rect 76579 7959 76637 7960
rect 76779 8000 76821 8009
rect 76779 7960 76780 8000
rect 76820 7960 76821 8000
rect 76779 7951 76821 7960
rect 76971 8000 77013 8009
rect 76971 7960 76972 8000
rect 77012 7960 77013 8000
rect 76971 7951 77013 7960
rect 77163 8000 77205 8009
rect 77163 7960 77164 8000
rect 77204 7960 77205 8000
rect 77163 7951 77205 7960
rect 77251 8000 77309 8001
rect 77251 7960 77260 8000
rect 77300 7960 77309 8000
rect 77251 7959 77309 7960
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 1219 7916 1277 7917
rect 1219 7876 1228 7916
rect 1268 7876 1277 7916
rect 1219 7875 1277 7876
rect 1611 7832 1653 7841
rect 1611 7792 1612 7832
rect 1652 7792 1653 7832
rect 1611 7783 1653 7792
rect 2763 7832 2805 7841
rect 2763 7792 2764 7832
rect 2804 7792 2805 7832
rect 2763 7783 2805 7792
rect 44427 7832 44469 7841
rect 44427 7792 44428 7832
rect 44468 7792 44469 7832
rect 44427 7783 44469 7792
rect 45867 7832 45909 7841
rect 45867 7792 45868 7832
rect 45908 7792 45909 7832
rect 45867 7783 45909 7792
rect 47019 7832 47061 7841
rect 47019 7792 47020 7832
rect 47060 7792 47061 7832
rect 47019 7783 47061 7792
rect 48643 7832 48701 7833
rect 48643 7792 48652 7832
rect 48692 7792 48701 7832
rect 48643 7791 48701 7792
rect 63051 7832 63093 7841
rect 63051 7792 63052 7832
rect 63092 7792 63093 7832
rect 63051 7783 63093 7792
rect 77739 7832 77781 7841
rect 77739 7792 77740 7832
rect 77780 7792 77781 7832
rect 77739 7783 77781 7792
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 1035 7748 1077 7757
rect 1035 7708 1036 7748
rect 1076 7708 1077 7748
rect 1035 7699 1077 7708
rect 4099 7748 4157 7749
rect 4099 7708 4108 7748
rect 4148 7708 4157 7748
rect 4099 7707 4157 7708
rect 7459 7748 7517 7749
rect 7459 7708 7468 7748
rect 7508 7708 7517 7748
rect 7459 7707 7517 7708
rect 47499 7748 47541 7757
rect 47499 7708 47500 7748
rect 47540 7708 47541 7748
rect 47499 7699 47541 7708
rect 49899 7748 49941 7757
rect 49899 7708 49900 7748
rect 49940 7708 49941 7748
rect 49899 7699 49941 7708
rect 58827 7748 58869 7757
rect 58827 7708 58828 7748
rect 58868 7708 58869 7748
rect 58827 7699 58869 7708
rect 60171 7748 60213 7757
rect 60171 7708 60172 7748
rect 60212 7708 60213 7748
rect 60171 7699 60213 7708
rect 63627 7748 63669 7757
rect 63627 7708 63628 7748
rect 63668 7708 63669 7748
rect 63627 7699 63669 7708
rect 65347 7748 65405 7749
rect 65347 7708 65356 7748
rect 65396 7708 65405 7748
rect 65347 7707 65405 7708
rect 68419 7748 68477 7749
rect 68419 7708 68428 7748
rect 68468 7708 68477 7748
rect 68419 7707 68477 7708
rect 71011 7748 71069 7749
rect 71011 7708 71020 7748
rect 71060 7708 71069 7748
rect 71011 7707 71069 7708
rect 76683 7748 76725 7757
rect 76683 7708 76684 7748
rect 76724 7708 76725 7748
rect 76683 7699 76725 7708
rect 576 7580 79584 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 79584 7580
rect 576 7516 79584 7540
rect 3907 7412 3965 7413
rect 3907 7372 3916 7412
rect 3956 7372 3965 7412
rect 3907 7371 3965 7372
rect 5067 7412 5109 7421
rect 5067 7372 5068 7412
rect 5108 7372 5109 7412
rect 5067 7363 5109 7372
rect 47779 7412 47837 7413
rect 47779 7372 47788 7412
rect 47828 7372 47837 7412
rect 47779 7371 47837 7372
rect 51139 7412 51197 7413
rect 51139 7372 51148 7412
rect 51188 7372 51197 7412
rect 51139 7371 51197 7372
rect 64579 7412 64637 7413
rect 64579 7372 64588 7412
rect 64628 7372 64637 7412
rect 64579 7371 64637 7372
rect 65355 7412 65397 7421
rect 65355 7372 65356 7412
rect 65396 7372 65397 7412
rect 65355 7363 65397 7372
rect 65931 7412 65973 7421
rect 65931 7372 65932 7412
rect 65972 7372 65973 7412
rect 65931 7363 65973 7372
rect 75531 7412 75573 7421
rect 75531 7372 75532 7412
rect 75572 7372 75573 7412
rect 75531 7363 75573 7372
rect 5547 7328 5589 7337
rect 5547 7288 5548 7328
rect 5588 7288 5589 7328
rect 5547 7279 5589 7288
rect 51915 7328 51957 7337
rect 51915 7288 51916 7328
rect 51956 7288 51957 7328
rect 51915 7279 51957 7288
rect 55083 7328 55125 7337
rect 55083 7288 55084 7328
rect 55124 7288 55125 7328
rect 55083 7279 55125 7288
rect 69387 7328 69429 7337
rect 69387 7288 69388 7328
rect 69428 7288 69429 7328
rect 69387 7279 69429 7288
rect 72459 7328 72501 7337
rect 72459 7288 72460 7328
rect 72500 7288 72501 7328
rect 72459 7279 72501 7288
rect 77835 7328 77877 7337
rect 77835 7288 77836 7328
rect 77876 7288 77877 7328
rect 77835 7279 77877 7288
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 54691 7244 54749 7245
rect 54691 7204 54700 7244
rect 54740 7204 54749 7244
rect 54691 7203 54749 7204
rect 76011 7171 76053 7180
rect 1891 7160 1949 7161
rect 1891 7120 1900 7160
rect 1940 7120 1949 7160
rect 1891 7119 1949 7120
rect 2755 7160 2813 7161
rect 2755 7120 2764 7160
rect 2804 7120 2813 7160
rect 2755 7119 2813 7120
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4387 7160 4445 7161
rect 4387 7120 4396 7160
rect 4436 7120 4445 7160
rect 4387 7119 4445 7120
rect 4963 7160 5021 7161
rect 4963 7120 4972 7160
rect 5012 7120 5021 7160
rect 4963 7119 5021 7120
rect 5163 7160 5205 7169
rect 5163 7120 5164 7160
rect 5204 7120 5205 7160
rect 5163 7111 5205 7120
rect 45387 7160 45429 7169
rect 45387 7120 45388 7160
rect 45428 7120 45429 7160
rect 45387 7111 45429 7120
rect 45763 7160 45821 7161
rect 45763 7120 45772 7160
rect 45812 7120 45821 7160
rect 45763 7119 45821 7120
rect 46627 7160 46685 7161
rect 46627 7120 46636 7160
rect 46676 7120 46685 7160
rect 46627 7119 46685 7120
rect 48747 7160 48789 7169
rect 48747 7120 48748 7160
rect 48788 7120 48789 7160
rect 48747 7111 48789 7120
rect 49123 7160 49181 7161
rect 49123 7120 49132 7160
rect 49172 7120 49181 7160
rect 49123 7119 49181 7120
rect 49987 7160 50045 7161
rect 49987 7120 49996 7160
rect 50036 7120 50045 7160
rect 49987 7119 50045 7120
rect 52779 7160 52821 7169
rect 52779 7120 52780 7160
rect 52820 7120 52821 7160
rect 52779 7111 52821 7120
rect 52971 7160 53013 7169
rect 52971 7120 52972 7160
rect 53012 7120 53013 7160
rect 52971 7111 53013 7120
rect 53059 7160 53117 7161
rect 53059 7120 53068 7160
rect 53108 7120 53117 7160
rect 53451 7160 53493 7169
rect 53059 7119 53117 7120
rect 53259 7118 53301 7127
rect 1515 7076 1557 7085
rect 1515 7036 1516 7076
rect 1556 7036 1557 7076
rect 1515 7027 1557 7036
rect 4299 7076 4341 7085
rect 4299 7036 4300 7076
rect 4340 7036 4341 7076
rect 4299 7027 4341 7036
rect 52875 7076 52917 7085
rect 52875 7036 52876 7076
rect 52916 7036 52917 7076
rect 53259 7078 53260 7118
rect 53300 7078 53301 7118
rect 53451 7120 53452 7160
rect 53492 7120 53493 7160
rect 53451 7111 53493 7120
rect 53539 7160 53597 7161
rect 53539 7120 53548 7160
rect 53588 7120 53597 7160
rect 53539 7119 53597 7120
rect 54307 7160 54365 7161
rect 54307 7120 54316 7160
rect 54356 7120 54365 7160
rect 54307 7119 54365 7120
rect 54507 7160 54549 7169
rect 54507 7120 54508 7160
rect 54548 7120 54549 7160
rect 54507 7111 54549 7120
rect 57187 7160 57245 7161
rect 57187 7120 57196 7160
rect 57236 7120 57245 7160
rect 57187 7119 57245 7120
rect 58051 7160 58109 7161
rect 58051 7120 58060 7160
rect 58100 7120 58109 7160
rect 58051 7119 58109 7120
rect 59683 7160 59741 7161
rect 59683 7120 59692 7160
rect 59732 7120 59741 7160
rect 59683 7119 59741 7120
rect 59979 7160 60021 7169
rect 59979 7120 59980 7160
rect 60020 7120 60021 7160
rect 59979 7111 60021 7120
rect 60547 7160 60605 7161
rect 60547 7120 60556 7160
rect 60596 7120 60605 7160
rect 60547 7119 60605 7120
rect 60651 7160 60693 7169
rect 60651 7120 60652 7160
rect 60692 7120 60693 7160
rect 60651 7111 60693 7120
rect 60843 7160 60885 7169
rect 60843 7120 60844 7160
rect 60884 7120 60885 7160
rect 60843 7111 60885 7120
rect 62187 7160 62229 7169
rect 62187 7120 62188 7160
rect 62228 7120 62229 7160
rect 62187 7111 62229 7120
rect 62563 7160 62621 7161
rect 62563 7120 62572 7160
rect 62612 7120 62621 7160
rect 62563 7119 62621 7120
rect 63427 7160 63485 7161
rect 63427 7120 63436 7160
rect 63476 7120 63485 7160
rect 63427 7119 63485 7120
rect 64779 7160 64821 7169
rect 64779 7120 64780 7160
rect 64820 7120 64821 7160
rect 64779 7111 64821 7120
rect 64971 7160 65013 7169
rect 64971 7120 64972 7160
rect 65012 7120 65013 7160
rect 64971 7111 65013 7120
rect 65059 7160 65117 7161
rect 65059 7120 65068 7160
rect 65108 7120 65117 7160
rect 65059 7119 65117 7120
rect 65251 7160 65309 7161
rect 65251 7120 65260 7160
rect 65300 7120 65309 7160
rect 65251 7119 65309 7120
rect 65451 7160 65493 7169
rect 65451 7120 65452 7160
rect 65492 7120 65493 7160
rect 65827 7161 65885 7162
rect 65827 7121 65836 7161
rect 65876 7121 65885 7161
rect 65827 7120 65885 7121
rect 66027 7160 66069 7169
rect 66027 7120 66028 7160
rect 66068 7120 66069 7160
rect 65451 7111 65493 7120
rect 66027 7111 66069 7120
rect 66211 7160 66269 7161
rect 66211 7120 66220 7160
rect 66260 7120 66269 7160
rect 66211 7119 66269 7120
rect 66411 7160 66453 7169
rect 66411 7120 66412 7160
rect 66452 7120 66453 7160
rect 66411 7111 66453 7120
rect 66595 7160 66653 7161
rect 66595 7120 66604 7160
rect 66644 7120 66653 7160
rect 66595 7119 66653 7120
rect 66795 7160 66837 7169
rect 66795 7120 66796 7160
rect 66836 7120 66837 7160
rect 66795 7111 66837 7120
rect 69579 7160 69621 7169
rect 69579 7120 69580 7160
rect 69620 7120 69621 7160
rect 69579 7111 69621 7120
rect 69675 7160 69717 7169
rect 69675 7120 69676 7160
rect 69716 7120 69717 7160
rect 69675 7111 69717 7120
rect 69771 7160 69813 7169
rect 69771 7120 69772 7160
rect 69812 7120 69813 7160
rect 69771 7111 69813 7120
rect 69867 7160 69909 7169
rect 69867 7120 69868 7160
rect 69908 7120 69909 7160
rect 69867 7111 69909 7120
rect 70059 7160 70101 7169
rect 70059 7120 70060 7160
rect 70100 7120 70101 7160
rect 70059 7111 70101 7120
rect 70251 7160 70293 7169
rect 70251 7120 70252 7160
rect 70292 7120 70293 7160
rect 70251 7111 70293 7120
rect 70339 7160 70397 7161
rect 70339 7120 70348 7160
rect 70388 7120 70397 7160
rect 70339 7119 70397 7120
rect 71691 7160 71733 7169
rect 71691 7120 71692 7160
rect 71732 7120 71733 7160
rect 71691 7111 71733 7120
rect 71883 7160 71925 7169
rect 71883 7120 71884 7160
rect 71924 7120 71925 7160
rect 71883 7111 71925 7120
rect 71971 7160 72029 7161
rect 71971 7120 71980 7160
rect 72020 7120 72029 7160
rect 71971 7119 72029 7120
rect 75531 7160 75573 7169
rect 75531 7120 75532 7160
rect 75572 7120 75573 7160
rect 75531 7111 75573 7120
rect 75723 7160 75765 7169
rect 75723 7120 75724 7160
rect 75764 7120 75765 7160
rect 75723 7111 75765 7120
rect 75811 7160 75869 7161
rect 75811 7120 75820 7160
rect 75860 7120 75869 7160
rect 76011 7131 76012 7171
rect 76052 7131 76053 7171
rect 76011 7122 76053 7131
rect 76203 7160 76245 7169
rect 75811 7119 75869 7120
rect 76203 7120 76204 7160
rect 76244 7120 76245 7160
rect 76203 7111 76245 7120
rect 76291 7160 76349 7161
rect 76291 7120 76300 7160
rect 76340 7120 76349 7160
rect 76291 7119 76349 7120
rect 76971 7160 77013 7169
rect 76971 7120 76972 7160
rect 77012 7120 77013 7160
rect 76971 7111 77013 7120
rect 77155 7160 77213 7161
rect 77155 7120 77164 7160
rect 77204 7120 77213 7160
rect 77155 7119 77213 7120
rect 77443 7160 77501 7161
rect 77443 7120 77452 7160
rect 77492 7120 77501 7160
rect 77443 7119 77501 7120
rect 77643 7160 77685 7169
rect 77643 7120 77644 7160
rect 77684 7120 77685 7160
rect 77643 7111 77685 7120
rect 53259 7069 53301 7078
rect 53355 7076 53397 7085
rect 52875 7027 52917 7036
rect 53355 7036 53356 7076
rect 53396 7036 53397 7076
rect 53355 7027 53397 7036
rect 54411 7076 54453 7085
rect 54411 7036 54412 7076
rect 54452 7036 54453 7076
rect 54411 7027 54453 7036
rect 56811 7076 56853 7085
rect 56811 7036 56812 7076
rect 56852 7036 56853 7076
rect 56811 7027 56853 7036
rect 60075 7076 60117 7085
rect 60075 7036 60076 7076
rect 60116 7036 60117 7076
rect 60075 7027 60117 7036
rect 60747 7076 60789 7085
rect 60747 7036 60748 7076
rect 60788 7036 60789 7076
rect 60747 7027 60789 7036
rect 64875 7076 64917 7085
rect 64875 7036 64876 7076
rect 64916 7036 64917 7076
rect 64875 7027 64917 7036
rect 66315 7076 66357 7085
rect 66315 7036 66316 7076
rect 66356 7036 66357 7076
rect 66315 7027 66357 7036
rect 66699 7076 66741 7085
rect 66699 7036 66700 7076
rect 66740 7036 66741 7076
rect 66699 7027 66741 7036
rect 76107 7076 76149 7085
rect 76107 7036 76108 7076
rect 76148 7036 76149 7076
rect 76107 7027 76149 7036
rect 77067 7076 77109 7085
rect 77067 7036 77068 7076
rect 77108 7036 77109 7076
rect 77067 7027 77109 7036
rect 77547 7076 77589 7085
rect 77547 7036 77548 7076
rect 77588 7036 77589 7076
rect 77547 7027 77589 7036
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 54891 6992 54933 7001
rect 54891 6952 54892 6992
rect 54932 6952 54933 6992
rect 54891 6943 54933 6952
rect 59203 6992 59261 6993
rect 59203 6952 59212 6992
rect 59252 6952 59261 6992
rect 70147 6992 70205 6993
rect 59203 6951 59261 6952
rect 60363 6950 60405 6959
rect 70147 6952 70156 6992
rect 70196 6952 70205 6992
rect 70147 6951 70205 6952
rect 71779 6992 71837 6993
rect 71779 6952 71788 6992
rect 71828 6952 71837 6992
rect 71779 6951 71837 6952
rect 60363 6910 60364 6950
rect 60404 6910 60405 6950
rect 60363 6901 60405 6910
rect 576 6824 79584 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 79584 6824
rect 576 6760 79584 6784
rect 2179 6656 2237 6657
rect 2179 6616 2188 6656
rect 2228 6616 2237 6656
rect 2179 6615 2237 6616
rect 7459 6656 7517 6657
rect 7459 6616 7468 6656
rect 7508 6616 7517 6656
rect 7459 6615 7517 6616
rect 47203 6656 47261 6657
rect 47203 6616 47212 6656
rect 47252 6616 47261 6656
rect 47203 6615 47261 6616
rect 53827 6656 53885 6657
rect 53827 6616 53836 6656
rect 53876 6616 53885 6656
rect 53827 6615 53885 6616
rect 56995 6656 57053 6657
rect 56995 6616 57004 6656
rect 57044 6616 57053 6656
rect 56995 6615 57053 6616
rect 68995 6656 69053 6657
rect 68995 6616 69004 6656
rect 69044 6616 69053 6656
rect 68995 6615 69053 6616
rect 74371 6656 74429 6657
rect 74371 6616 74380 6656
rect 74420 6616 74429 6656
rect 74371 6615 74429 6616
rect 79459 6656 79517 6657
rect 79459 6616 79468 6656
rect 79508 6616 79517 6656
rect 79459 6615 79517 6616
rect 54219 6572 54261 6581
rect 54219 6532 54220 6572
rect 54260 6532 54261 6572
rect 54219 6523 54261 6532
rect 54603 6572 54645 6581
rect 54603 6532 54604 6572
rect 54644 6532 54645 6572
rect 54603 6523 54645 6532
rect 66027 6572 66069 6581
rect 66027 6532 66028 6572
rect 66068 6532 66069 6572
rect 66027 6523 66069 6532
rect 71979 6572 72021 6581
rect 71979 6532 71980 6572
rect 72020 6532 72021 6572
rect 71979 6523 72021 6532
rect 2091 6488 2133 6497
rect 2091 6448 2092 6488
rect 2132 6448 2133 6488
rect 2091 6439 2133 6448
rect 2283 6488 2325 6497
rect 2283 6448 2284 6488
rect 2324 6448 2325 6488
rect 2283 6439 2325 6448
rect 2371 6488 2429 6489
rect 2371 6448 2380 6488
rect 2420 6448 2429 6488
rect 2371 6447 2429 6448
rect 2571 6488 2613 6497
rect 2571 6448 2572 6488
rect 2612 6448 2613 6488
rect 2571 6439 2613 6448
rect 2763 6488 2805 6497
rect 2763 6448 2764 6488
rect 2804 6448 2805 6488
rect 4107 6488 4149 6497
rect 2763 6439 2805 6448
rect 2861 6469 2919 6470
rect 2861 6429 2870 6469
rect 2910 6429 2919 6469
rect 4107 6448 4108 6488
rect 4148 6448 4149 6488
rect 4107 6439 4149 6448
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 4483 6488 4541 6489
rect 4483 6448 4492 6488
rect 4532 6448 4541 6488
rect 4483 6447 4541 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5443 6488 5501 6489
rect 5443 6448 5452 6488
rect 5492 6448 5501 6488
rect 5443 6447 5501 6448
rect 6307 6488 6365 6489
rect 6307 6448 6316 6488
rect 6356 6448 6365 6488
rect 6307 6447 6365 6448
rect 47307 6488 47349 6497
rect 47307 6448 47308 6488
rect 47348 6448 47349 6488
rect 47307 6439 47349 6448
rect 47403 6488 47445 6497
rect 47403 6448 47404 6488
rect 47444 6448 47445 6488
rect 47403 6439 47445 6448
rect 47499 6488 47541 6497
rect 47499 6448 47500 6488
rect 47540 6448 47541 6488
rect 47499 6439 47541 6448
rect 47691 6488 47733 6497
rect 47691 6448 47692 6488
rect 47732 6448 47733 6488
rect 47691 6439 47733 6448
rect 47883 6488 47925 6497
rect 47883 6448 47884 6488
rect 47924 6448 47925 6488
rect 47883 6439 47925 6448
rect 47971 6488 48029 6489
rect 47971 6448 47980 6488
rect 48020 6448 48029 6488
rect 47971 6447 48029 6448
rect 48355 6488 48413 6489
rect 48355 6448 48364 6488
rect 48404 6448 48413 6488
rect 48355 6447 48413 6448
rect 48555 6488 48597 6497
rect 48555 6448 48556 6488
rect 48596 6448 48597 6488
rect 48555 6439 48597 6448
rect 48843 6488 48885 6497
rect 48843 6448 48844 6488
rect 48884 6448 48885 6488
rect 48843 6439 48885 6448
rect 49219 6488 49277 6489
rect 49219 6448 49228 6488
rect 49268 6448 49277 6488
rect 49219 6447 49277 6448
rect 50083 6488 50141 6489
rect 50083 6448 50092 6488
rect 50132 6448 50141 6488
rect 50083 6447 50141 6448
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51811 6488 51869 6489
rect 51811 6448 51820 6488
rect 51860 6448 51869 6488
rect 51811 6447 51869 6448
rect 52675 6488 52733 6489
rect 52675 6448 52684 6488
rect 52724 6448 52733 6488
rect 52675 6447 52733 6448
rect 54123 6488 54165 6497
rect 54123 6448 54124 6488
rect 54164 6448 54165 6488
rect 54123 6439 54165 6448
rect 54315 6488 54357 6497
rect 54315 6448 54316 6488
rect 54356 6448 54357 6488
rect 54315 6439 54357 6448
rect 54403 6488 54461 6489
rect 54403 6448 54412 6488
rect 54452 6448 54461 6488
rect 54403 6447 54461 6448
rect 54979 6488 55037 6489
rect 54979 6448 54988 6488
rect 55028 6448 55037 6488
rect 54979 6447 55037 6448
rect 55843 6488 55901 6489
rect 55843 6448 55852 6488
rect 55892 6448 55901 6488
rect 55843 6447 55901 6448
rect 58059 6488 58101 6497
rect 58059 6448 58060 6488
rect 58100 6448 58101 6488
rect 58059 6439 58101 6448
rect 58251 6488 58293 6497
rect 58251 6448 58252 6488
rect 58292 6448 58293 6488
rect 58251 6439 58293 6448
rect 58339 6488 58397 6489
rect 58339 6448 58348 6488
rect 58388 6448 58397 6488
rect 58339 6447 58397 6448
rect 58539 6488 58581 6497
rect 58539 6448 58540 6488
rect 58580 6448 58581 6488
rect 58539 6439 58581 6448
rect 58635 6488 58677 6497
rect 58635 6448 58636 6488
rect 58676 6448 58677 6488
rect 58635 6439 58677 6448
rect 58731 6488 58773 6497
rect 58731 6448 58732 6488
rect 58772 6448 58773 6488
rect 58731 6439 58773 6448
rect 58827 6488 58869 6497
rect 58827 6448 58828 6488
rect 58868 6448 58869 6488
rect 58827 6439 58869 6448
rect 59203 6488 59261 6489
rect 59203 6448 59212 6488
rect 59252 6448 59261 6488
rect 59203 6447 59261 6448
rect 59307 6488 59349 6497
rect 59307 6448 59308 6488
rect 59348 6448 59349 6488
rect 59307 6439 59349 6448
rect 59499 6488 59541 6497
rect 59499 6448 59500 6488
rect 59540 6448 59541 6488
rect 59499 6439 59541 6448
rect 60163 6488 60221 6489
rect 60163 6448 60172 6488
rect 60212 6448 60221 6488
rect 60163 6447 60221 6448
rect 60363 6488 60405 6497
rect 60363 6448 60364 6488
rect 60404 6448 60405 6488
rect 60363 6439 60405 6448
rect 61035 6488 61077 6497
rect 61035 6448 61036 6488
rect 61076 6448 61077 6488
rect 61035 6439 61077 6448
rect 61227 6488 61269 6497
rect 61227 6448 61228 6488
rect 61268 6448 61269 6488
rect 61227 6439 61269 6448
rect 61315 6488 61373 6489
rect 61315 6448 61324 6488
rect 61364 6448 61373 6488
rect 61315 6447 61373 6448
rect 65635 6488 65693 6489
rect 65635 6448 65644 6488
rect 65684 6448 65693 6488
rect 65635 6447 65693 6448
rect 65931 6488 65973 6497
rect 65931 6448 65932 6488
rect 65972 6448 65973 6488
rect 65931 6439 65973 6448
rect 66603 6488 66645 6497
rect 66603 6448 66604 6488
rect 66644 6448 66645 6488
rect 66603 6439 66645 6448
rect 66979 6488 67037 6489
rect 66979 6448 66988 6488
rect 67028 6448 67037 6488
rect 66979 6447 67037 6448
rect 67843 6488 67901 6489
rect 67843 6448 67852 6488
rect 67892 6448 67901 6488
rect 67843 6447 67901 6448
rect 69195 6488 69237 6497
rect 69195 6448 69196 6488
rect 69236 6448 69237 6488
rect 69195 6439 69237 6448
rect 69571 6488 69629 6489
rect 69571 6448 69580 6488
rect 69620 6448 69629 6488
rect 69571 6447 69629 6448
rect 70435 6488 70493 6489
rect 70435 6448 70444 6488
rect 70484 6448 70493 6488
rect 70435 6447 70493 6448
rect 72355 6488 72413 6489
rect 72355 6448 72364 6488
rect 72404 6448 72413 6488
rect 72355 6447 72413 6448
rect 73219 6488 73277 6489
rect 73219 6448 73228 6488
rect 73268 6448 73277 6488
rect 73219 6447 73277 6448
rect 75627 6488 75669 6497
rect 75627 6448 75628 6488
rect 75668 6448 75669 6488
rect 75627 6439 75669 6448
rect 75723 6488 75765 6497
rect 75723 6448 75724 6488
rect 75764 6448 75765 6488
rect 75723 6439 75765 6448
rect 75819 6488 75861 6497
rect 75819 6448 75820 6488
rect 75860 6448 75861 6488
rect 75819 6439 75861 6448
rect 75915 6488 75957 6497
rect 75915 6448 75916 6488
rect 75956 6448 75957 6488
rect 75915 6439 75957 6448
rect 76195 6488 76253 6489
rect 76195 6448 76204 6488
rect 76244 6448 76253 6488
rect 76195 6447 76253 6448
rect 76491 6488 76533 6497
rect 76491 6448 76492 6488
rect 76532 6448 76533 6488
rect 76491 6439 76533 6448
rect 76587 6488 76629 6497
rect 76587 6448 76588 6488
rect 76628 6448 76629 6488
rect 76587 6439 76629 6448
rect 77067 6488 77109 6497
rect 77067 6448 77068 6488
rect 77108 6448 77109 6488
rect 77067 6439 77109 6448
rect 77443 6488 77501 6489
rect 77443 6448 77452 6488
rect 77492 6448 77501 6488
rect 77443 6447 77501 6448
rect 78307 6488 78365 6489
rect 78307 6448 78316 6488
rect 78356 6448 78365 6488
rect 78307 6447 78365 6448
rect 2861 6428 2919 6429
rect 1707 6320 1749 6329
rect 1707 6280 1708 6320
rect 1748 6280 1749 6320
rect 1707 6271 1749 6280
rect 2571 6320 2613 6329
rect 2571 6280 2572 6320
rect 2612 6280 2613 6320
rect 2571 6271 2613 6280
rect 57291 6320 57333 6329
rect 57291 6280 57292 6320
rect 57332 6280 57333 6320
rect 57291 6271 57333 6280
rect 58059 6320 58101 6329
rect 58059 6280 58060 6320
rect 58100 6280 58101 6320
rect 58059 6271 58101 6280
rect 60267 6320 60309 6329
rect 60267 6280 60268 6320
rect 60308 6280 60309 6320
rect 60267 6271 60309 6280
rect 61707 6320 61749 6329
rect 61707 6280 61708 6320
rect 61748 6280 61749 6320
rect 61707 6271 61749 6280
rect 63435 6320 63477 6329
rect 63435 6280 63436 6320
rect 63476 6280 63477 6320
rect 63435 6271 63477 6280
rect 66307 6320 66365 6321
rect 66307 6280 66316 6320
rect 66356 6280 66365 6320
rect 66307 6279 66365 6280
rect 74763 6320 74805 6329
rect 74763 6280 74764 6320
rect 74804 6280 74805 6320
rect 74763 6271 74805 6280
rect 76867 6320 76925 6321
rect 76867 6280 76876 6320
rect 76916 6280 76925 6320
rect 76867 6279 76925 6280
rect 3811 6236 3869 6237
rect 3811 6196 3820 6236
rect 3860 6196 3869 6236
rect 3811 6195 3869 6196
rect 47691 6236 47733 6245
rect 47691 6196 47692 6236
rect 47732 6196 47733 6236
rect 47691 6187 47733 6196
rect 48459 6236 48501 6245
rect 48459 6196 48460 6236
rect 48500 6196 48501 6236
rect 48459 6187 48501 6196
rect 51235 6236 51293 6237
rect 51235 6196 51244 6236
rect 51284 6196 51293 6236
rect 51235 6195 51293 6196
rect 53827 6236 53885 6237
rect 53827 6196 53836 6236
rect 53876 6196 53885 6236
rect 53827 6195 53885 6196
rect 56995 6236 57053 6237
rect 56995 6196 57004 6236
rect 57044 6196 57053 6236
rect 56995 6195 57053 6196
rect 59499 6236 59541 6245
rect 59499 6196 59500 6236
rect 59540 6196 59541 6236
rect 59499 6187 59541 6196
rect 61035 6236 61077 6245
rect 61035 6196 61036 6236
rect 61076 6196 61077 6236
rect 61035 6187 61077 6196
rect 71587 6236 71645 6237
rect 71587 6196 71596 6236
rect 71636 6196 71645 6236
rect 71587 6195 71645 6196
rect 74371 6236 74429 6237
rect 74371 6196 74380 6236
rect 74420 6196 74429 6236
rect 74371 6195 74429 6196
rect 576 6068 79584 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 79584 6068
rect 576 6004 79584 6028
rect 6315 5900 6357 5909
rect 6315 5860 6316 5900
rect 6356 5860 6357 5900
rect 6315 5851 6357 5860
rect 48739 5900 48797 5901
rect 48739 5860 48748 5900
rect 48788 5860 48797 5900
rect 48739 5859 48797 5860
rect 48939 5900 48981 5909
rect 48939 5860 48940 5900
rect 48980 5860 48981 5900
rect 48939 5851 48981 5860
rect 54499 5900 54557 5901
rect 54499 5860 54508 5900
rect 54548 5860 54557 5900
rect 54499 5859 54557 5860
rect 66315 5900 66357 5909
rect 66315 5860 66316 5900
rect 66356 5860 66357 5900
rect 66315 5851 66357 5860
rect 69771 5900 69813 5909
rect 69771 5860 69772 5900
rect 69812 5860 69813 5900
rect 69771 5851 69813 5860
rect 72651 5900 72693 5909
rect 72651 5860 72652 5900
rect 72692 5860 72693 5900
rect 72651 5851 72693 5860
rect 73603 5900 73661 5901
rect 73603 5860 73612 5900
rect 73652 5860 73661 5900
rect 73603 5859 73661 5860
rect 77163 5900 77205 5909
rect 77163 5860 77164 5900
rect 77204 5860 77205 5900
rect 77163 5851 77205 5860
rect 46155 5816 46197 5825
rect 46155 5776 46156 5816
rect 46196 5776 46197 5816
rect 46155 5767 46197 5776
rect 49419 5816 49461 5825
rect 49419 5776 49420 5816
rect 49460 5776 49461 5816
rect 49419 5767 49461 5776
rect 56619 5816 56661 5825
rect 56619 5776 56620 5816
rect 56660 5776 56661 5816
rect 56619 5767 56661 5776
rect 59691 5816 59733 5825
rect 59691 5776 59692 5816
rect 59732 5776 59733 5816
rect 59691 5767 59733 5776
rect 61027 5816 61085 5817
rect 61027 5776 61036 5816
rect 61076 5776 61085 5816
rect 61027 5775 61085 5776
rect 67179 5816 67221 5825
rect 67179 5776 67180 5816
rect 67220 5776 67221 5816
rect 67179 5767 67221 5776
rect 71971 5816 72029 5817
rect 71971 5776 71980 5816
rect 72020 5776 72029 5816
rect 71971 5775 72029 5776
rect 1027 5732 1085 5733
rect 1027 5692 1036 5732
rect 1076 5692 1085 5732
rect 1027 5691 1085 5692
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 54795 5732 54837 5741
rect 54795 5692 54796 5732
rect 54836 5692 54837 5732
rect 54795 5683 54837 5692
rect 1603 5648 1661 5649
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1603 5607 1661 5608
rect 2467 5648 2525 5649
rect 2467 5608 2476 5648
rect 2516 5608 2525 5648
rect 2467 5607 2525 5608
rect 5739 5648 5781 5657
rect 5739 5608 5740 5648
rect 5780 5608 5781 5648
rect 5739 5599 5781 5608
rect 6019 5648 6077 5649
rect 6019 5608 6028 5648
rect 6068 5608 6077 5648
rect 6019 5607 6077 5608
rect 6123 5648 6165 5657
rect 6123 5608 6124 5648
rect 6164 5608 6165 5648
rect 6123 5599 6165 5608
rect 6315 5648 6357 5657
rect 6315 5608 6316 5648
rect 6356 5608 6357 5648
rect 6315 5599 6357 5608
rect 47211 5648 47253 5657
rect 47211 5608 47212 5648
rect 47252 5608 47253 5648
rect 47211 5599 47253 5608
rect 47403 5648 47445 5657
rect 47403 5608 47404 5648
rect 47444 5608 47445 5648
rect 47403 5599 47445 5608
rect 47491 5648 47549 5649
rect 47491 5608 47500 5648
rect 47540 5608 47549 5648
rect 47491 5607 47549 5608
rect 48067 5648 48125 5649
rect 48067 5608 48076 5648
rect 48116 5608 48125 5648
rect 48067 5607 48125 5608
rect 48363 5648 48405 5657
rect 48363 5608 48364 5648
rect 48404 5608 48405 5648
rect 48363 5599 48405 5608
rect 48939 5648 48981 5657
rect 48939 5608 48940 5648
rect 48980 5608 48981 5648
rect 48939 5599 48981 5608
rect 49131 5648 49173 5657
rect 49131 5608 49132 5648
rect 49172 5608 49173 5648
rect 49131 5599 49173 5608
rect 49219 5648 49277 5649
rect 49219 5608 49228 5648
rect 49268 5608 49277 5648
rect 49219 5607 49277 5608
rect 52195 5648 52253 5649
rect 52195 5608 52204 5648
rect 52244 5608 52253 5648
rect 52195 5607 52253 5608
rect 52299 5648 52341 5657
rect 52299 5608 52300 5648
rect 52340 5608 52341 5648
rect 52299 5599 52341 5608
rect 52491 5648 52533 5657
rect 52491 5608 52492 5648
rect 52532 5608 52533 5648
rect 52491 5599 52533 5608
rect 52779 5648 52821 5657
rect 52779 5608 52780 5648
rect 52820 5608 52821 5648
rect 52779 5599 52821 5608
rect 52875 5648 52917 5657
rect 52875 5608 52876 5648
rect 52916 5608 52917 5648
rect 52875 5599 52917 5608
rect 52971 5648 53013 5657
rect 52971 5608 52972 5648
rect 53012 5608 53013 5648
rect 52971 5599 53013 5608
rect 53827 5648 53885 5649
rect 53827 5608 53836 5648
rect 53876 5608 53885 5648
rect 53827 5607 53885 5608
rect 54123 5648 54165 5657
rect 54123 5608 54124 5648
rect 54164 5608 54165 5648
rect 54123 5599 54165 5608
rect 54219 5648 54261 5657
rect 54219 5608 54220 5648
rect 54260 5608 54261 5648
rect 54219 5599 54261 5608
rect 54699 5648 54741 5657
rect 54699 5608 54700 5648
rect 54740 5608 54741 5648
rect 54699 5599 54741 5608
rect 54883 5648 54941 5649
rect 54883 5608 54892 5648
rect 54932 5608 54941 5648
rect 54883 5607 54941 5608
rect 56227 5648 56285 5649
rect 56227 5608 56236 5648
rect 56276 5608 56285 5648
rect 56227 5607 56285 5608
rect 56427 5648 56469 5657
rect 56427 5608 56428 5648
rect 56468 5608 56469 5648
rect 56427 5599 56469 5608
rect 59211 5648 59253 5657
rect 59211 5608 59212 5648
rect 59252 5608 59253 5648
rect 59211 5599 59253 5608
rect 59403 5648 59445 5657
rect 59403 5608 59404 5648
rect 59444 5608 59445 5648
rect 59403 5599 59445 5608
rect 59491 5648 59549 5649
rect 59491 5608 59500 5648
rect 59540 5608 59549 5648
rect 59491 5607 59549 5608
rect 60355 5648 60413 5649
rect 60355 5608 60364 5648
rect 60404 5608 60413 5648
rect 60355 5607 60413 5608
rect 60651 5648 60693 5657
rect 60651 5608 60652 5648
rect 60692 5608 60693 5648
rect 60651 5599 60693 5608
rect 61227 5648 61269 5657
rect 61227 5608 61228 5648
rect 61268 5608 61269 5648
rect 61227 5599 61269 5608
rect 61603 5648 61661 5649
rect 61603 5608 61612 5648
rect 61652 5608 61661 5648
rect 61603 5607 61661 5608
rect 62467 5648 62525 5649
rect 62467 5608 62476 5648
rect 62516 5608 62525 5648
rect 62467 5607 62525 5608
rect 64587 5648 64629 5657
rect 64587 5608 64588 5648
rect 64628 5608 64629 5648
rect 64587 5599 64629 5608
rect 64779 5648 64821 5657
rect 64779 5608 64780 5648
rect 64820 5608 64821 5648
rect 64779 5599 64821 5608
rect 64867 5648 64925 5649
rect 64867 5608 64876 5648
rect 64916 5608 64925 5648
rect 64867 5607 64925 5608
rect 65067 5648 65109 5657
rect 65067 5608 65068 5648
rect 65108 5608 65109 5648
rect 65067 5599 65109 5608
rect 65163 5648 65205 5657
rect 65163 5608 65164 5648
rect 65204 5608 65205 5648
rect 65163 5599 65205 5608
rect 65259 5648 65301 5657
rect 65259 5608 65260 5648
rect 65300 5608 65301 5648
rect 65259 5599 65301 5608
rect 65355 5648 65397 5657
rect 65355 5608 65356 5648
rect 65396 5608 65397 5648
rect 66507 5648 66549 5657
rect 65355 5599 65397 5608
rect 66315 5606 66357 5615
rect 1227 5564 1269 5573
rect 1227 5524 1228 5564
rect 1268 5524 1269 5564
rect 1227 5515 1269 5524
rect 48459 5564 48501 5573
rect 48459 5524 48460 5564
rect 48500 5524 48501 5564
rect 48459 5515 48501 5524
rect 52395 5564 52437 5573
rect 52395 5524 52396 5564
rect 52436 5524 52437 5564
rect 52395 5515 52437 5524
rect 52683 5564 52725 5573
rect 52683 5524 52684 5564
rect 52724 5524 52725 5564
rect 52683 5515 52725 5524
rect 56331 5564 56373 5573
rect 56331 5524 56332 5564
rect 56372 5524 56373 5564
rect 56331 5515 56373 5524
rect 60747 5564 60789 5573
rect 60747 5524 60748 5564
rect 60788 5524 60789 5564
rect 66315 5566 66316 5606
rect 66356 5566 66357 5606
rect 66507 5608 66508 5648
rect 66548 5608 66549 5648
rect 66507 5599 66549 5608
rect 66595 5648 66653 5649
rect 66595 5608 66604 5648
rect 66644 5608 66653 5648
rect 69387 5648 69429 5657
rect 66595 5607 66653 5608
rect 69291 5627 69333 5636
rect 69291 5587 69292 5627
rect 69332 5587 69333 5627
rect 69387 5608 69388 5648
rect 69428 5608 69429 5648
rect 69387 5599 69429 5608
rect 69483 5648 69525 5657
rect 69483 5608 69484 5648
rect 69524 5608 69525 5648
rect 69483 5599 69525 5608
rect 69579 5648 69621 5657
rect 69579 5608 69580 5648
rect 69620 5608 69621 5648
rect 69579 5599 69621 5608
rect 69771 5648 69813 5657
rect 69771 5608 69772 5648
rect 69812 5608 69813 5648
rect 69771 5599 69813 5608
rect 69963 5648 70005 5657
rect 69963 5608 69964 5648
rect 70004 5608 70005 5648
rect 69963 5599 70005 5608
rect 70051 5648 70109 5649
rect 70051 5608 70060 5648
rect 70100 5608 70109 5648
rect 70051 5607 70109 5608
rect 71299 5648 71357 5649
rect 71299 5608 71308 5648
rect 71348 5608 71357 5648
rect 71299 5607 71357 5608
rect 71595 5648 71637 5657
rect 71595 5608 71596 5648
rect 71636 5608 71637 5648
rect 71595 5599 71637 5608
rect 71691 5648 71733 5657
rect 71691 5608 71692 5648
rect 71732 5608 71733 5648
rect 71691 5599 71733 5608
rect 72171 5648 72213 5657
rect 72171 5608 72172 5648
rect 72212 5608 72213 5648
rect 72171 5599 72213 5608
rect 72355 5648 72413 5649
rect 72355 5608 72364 5648
rect 72404 5608 72413 5648
rect 72355 5607 72413 5608
rect 72547 5648 72605 5649
rect 72547 5608 72556 5648
rect 72596 5608 72605 5648
rect 72547 5607 72605 5608
rect 72747 5648 72789 5657
rect 72747 5608 72748 5648
rect 72788 5608 72789 5648
rect 72747 5599 72789 5608
rect 74755 5648 74813 5649
rect 74755 5608 74764 5648
rect 74804 5608 74813 5648
rect 74755 5607 74813 5608
rect 75619 5648 75677 5649
rect 75619 5608 75628 5648
rect 75668 5608 75677 5648
rect 75619 5607 75677 5608
rect 76203 5648 76245 5657
rect 76203 5608 76204 5648
rect 76244 5608 76245 5648
rect 76203 5599 76245 5608
rect 76395 5648 76437 5657
rect 76395 5608 76396 5648
rect 76436 5608 76437 5648
rect 76395 5599 76437 5608
rect 76483 5648 76541 5649
rect 76483 5608 76492 5648
rect 76532 5608 76541 5648
rect 76483 5607 76541 5608
rect 77163 5648 77205 5657
rect 77163 5608 77164 5648
rect 77204 5608 77205 5648
rect 77163 5599 77205 5608
rect 77355 5648 77397 5657
rect 77355 5608 77356 5648
rect 77396 5608 77397 5648
rect 77355 5599 77397 5608
rect 77443 5648 77501 5649
rect 77443 5608 77452 5648
rect 77492 5608 77501 5648
rect 77443 5607 77501 5608
rect 69291 5578 69333 5587
rect 66315 5557 66357 5566
rect 72267 5564 72309 5573
rect 60747 5515 60789 5524
rect 72267 5524 72268 5564
rect 72308 5524 72309 5564
rect 72267 5515 72309 5524
rect 76011 5564 76053 5573
rect 76011 5524 76012 5564
rect 76052 5524 76053 5564
rect 76011 5515 76053 5524
rect 843 5480 885 5489
rect 843 5440 844 5480
rect 884 5440 885 5480
rect 843 5431 885 5440
rect 47299 5480 47357 5481
rect 47299 5440 47308 5480
rect 47348 5440 47357 5480
rect 47299 5439 47357 5440
rect 59299 5480 59357 5481
rect 59299 5440 59308 5480
rect 59348 5440 59357 5480
rect 59299 5439 59357 5440
rect 63619 5480 63677 5481
rect 63619 5440 63628 5480
rect 63668 5440 63677 5480
rect 63619 5439 63677 5440
rect 64675 5480 64733 5481
rect 64675 5440 64684 5480
rect 64724 5440 64733 5480
rect 64675 5439 64733 5440
rect 76291 5480 76349 5481
rect 76291 5440 76300 5480
rect 76340 5440 76349 5480
rect 76291 5439 76349 5440
rect 576 5312 79584 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 79584 5312
rect 576 5248 79584 5272
rect 651 5144 693 5153
rect 651 5104 652 5144
rect 692 5104 693 5144
rect 651 5095 693 5104
rect 2179 5144 2237 5145
rect 2179 5104 2188 5144
rect 2228 5104 2237 5144
rect 2179 5103 2237 5104
rect 52195 5144 52253 5145
rect 52195 5104 52204 5144
rect 52244 5104 52253 5144
rect 52195 5103 52253 5104
rect 55747 5144 55805 5145
rect 55747 5104 55756 5144
rect 55796 5104 55805 5144
rect 55747 5103 55805 5104
rect 65347 5144 65405 5145
rect 65347 5104 65356 5144
rect 65396 5104 65405 5144
rect 65347 5103 65405 5104
rect 65635 5144 65693 5145
rect 65635 5104 65644 5144
rect 65684 5104 65693 5144
rect 65635 5103 65693 5104
rect 76099 5144 76157 5145
rect 76099 5104 76108 5144
rect 76148 5104 76157 5144
rect 76099 5103 76157 5104
rect 3531 5060 3573 5069
rect 3531 5020 3532 5060
rect 3572 5020 3573 5060
rect 3531 5011 3573 5020
rect 3915 5060 3957 5069
rect 3915 5020 3916 5060
rect 3956 5020 3957 5060
rect 3915 5011 3957 5020
rect 4291 5060 4349 5061
rect 4291 5020 4300 5060
rect 4340 5020 4349 5060
rect 4291 5019 4349 5020
rect 45675 5060 45717 5069
rect 45675 5020 45676 5060
rect 45716 5020 45717 5060
rect 45675 5011 45717 5020
rect 48555 5060 48597 5069
rect 48555 5020 48556 5060
rect 48596 5020 48597 5060
rect 48555 5011 48597 5020
rect 52587 5060 52629 5069
rect 52587 5020 52588 5060
rect 52628 5020 52629 5060
rect 52587 5011 52629 5020
rect 56139 5060 56181 5069
rect 56139 5020 56140 5060
rect 56180 5020 56181 5060
rect 56139 5011 56181 5020
rect 58827 5060 58869 5069
rect 58827 5020 58828 5060
rect 58868 5020 58869 5060
rect 58827 5011 58869 5020
rect 61899 5060 61941 5069
rect 61899 5020 61900 5060
rect 61940 5020 61941 5060
rect 61899 5011 61941 5020
rect 62955 5060 62997 5069
rect 62955 5020 62956 5060
rect 62996 5020 62997 5060
rect 62955 5011 62997 5020
rect 1611 4976 1653 4985
rect 1611 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 1707 4976 1749 4985
rect 1707 4936 1708 4976
rect 1748 4936 1749 4976
rect 1707 4927 1749 4936
rect 1803 4976 1845 4985
rect 1803 4936 1804 4976
rect 1844 4936 1845 4976
rect 1803 4927 1845 4936
rect 1899 4976 1941 4985
rect 1899 4936 1900 4976
rect 1940 4936 1941 4976
rect 1899 4927 1941 4936
rect 2091 4976 2133 4985
rect 2091 4936 2092 4976
rect 2132 4936 2133 4976
rect 2091 4927 2133 4936
rect 2283 4976 2325 4985
rect 2283 4936 2284 4976
rect 2324 4936 2325 4976
rect 2283 4927 2325 4936
rect 2371 4976 2429 4977
rect 2371 4936 2380 4976
rect 2420 4936 2429 4976
rect 2371 4935 2429 4936
rect 3427 4976 3485 4977
rect 3427 4936 3436 4976
rect 3476 4936 3485 4976
rect 3427 4935 3485 4936
rect 3627 4976 3669 4985
rect 3627 4936 3628 4976
rect 3668 4936 3669 4976
rect 3627 4927 3669 4936
rect 3819 4976 3861 4985
rect 3819 4936 3820 4976
rect 3860 4936 3861 4976
rect 3819 4927 3861 4936
rect 4003 4976 4061 4977
rect 4003 4936 4012 4976
rect 4052 4936 4061 4976
rect 4003 4935 4061 4936
rect 5155 4976 5213 4977
rect 5155 4936 5164 4976
rect 5204 4936 5213 4976
rect 5155 4935 5213 4936
rect 46051 4976 46109 4977
rect 46051 4936 46060 4976
rect 46100 4936 46109 4976
rect 46051 4935 46109 4936
rect 46915 4976 46973 4977
rect 46915 4936 46924 4976
rect 46964 4936 46973 4976
rect 46915 4935 46973 4936
rect 48459 4976 48501 4985
rect 48459 4936 48460 4976
rect 48500 4936 48501 4976
rect 48459 4927 48501 4936
rect 48643 4976 48701 4977
rect 48643 4936 48652 4976
rect 48692 4936 48701 4976
rect 48643 4935 48701 4936
rect 48835 4976 48893 4977
rect 48835 4936 48844 4976
rect 48884 4936 48893 4976
rect 48835 4935 48893 4936
rect 48939 4976 48981 4985
rect 48939 4936 48940 4976
rect 48980 4936 48981 4976
rect 48939 4927 48981 4936
rect 49131 4976 49173 4985
rect 49131 4936 49132 4976
rect 49172 4936 49173 4976
rect 49131 4927 49173 4936
rect 51531 4976 51573 4985
rect 51531 4936 51532 4976
rect 51572 4936 51573 4976
rect 51531 4927 51573 4936
rect 51723 4976 51765 4985
rect 51723 4936 51724 4976
rect 51764 4936 51765 4976
rect 51723 4927 51765 4936
rect 51811 4976 51869 4977
rect 51811 4936 51820 4976
rect 51860 4936 51869 4976
rect 51811 4935 51869 4936
rect 52003 4976 52061 4977
rect 52003 4936 52012 4976
rect 52052 4936 52061 4976
rect 52003 4935 52061 4936
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 52299 4976 52341 4985
rect 52299 4936 52300 4976
rect 52340 4936 52341 4976
rect 52299 4927 52341 4936
rect 52483 4976 52541 4977
rect 52483 4936 52492 4976
rect 52532 4936 52541 4976
rect 52483 4935 52541 4936
rect 52683 4976 52725 4985
rect 52683 4936 52684 4976
rect 52724 4936 52725 4976
rect 52683 4927 52725 4936
rect 55659 4976 55701 4985
rect 55659 4936 55660 4976
rect 55700 4936 55701 4976
rect 55659 4927 55701 4936
rect 55851 4976 55893 4985
rect 55851 4936 55852 4976
rect 55892 4936 55893 4976
rect 55851 4927 55893 4936
rect 55939 4976 55997 4977
rect 55939 4936 55948 4976
rect 55988 4936 55997 4976
rect 55939 4935 55997 4936
rect 56515 4976 56573 4977
rect 56515 4936 56524 4976
rect 56564 4936 56573 4976
rect 56515 4935 56573 4936
rect 57379 4976 57437 4977
rect 57379 4936 57388 4976
rect 57428 4936 57437 4976
rect 57379 4935 57437 4936
rect 59203 4976 59261 4977
rect 59203 4936 59212 4976
rect 59252 4936 59261 4976
rect 59203 4935 59261 4936
rect 60067 4976 60125 4977
rect 60067 4936 60076 4976
rect 60116 4936 60125 4976
rect 60067 4935 60125 4936
rect 61419 4976 61461 4985
rect 61419 4936 61420 4976
rect 61460 4936 61461 4976
rect 61419 4927 61461 4936
rect 61603 4976 61661 4977
rect 61603 4936 61612 4976
rect 61652 4936 61661 4976
rect 61603 4935 61661 4936
rect 61795 4976 61853 4977
rect 61795 4936 61804 4976
rect 61844 4936 61853 4976
rect 61795 4935 61853 4936
rect 61995 4976 62037 4985
rect 61995 4936 61996 4976
rect 62036 4936 62037 4976
rect 61995 4927 62037 4936
rect 63331 4976 63389 4977
rect 63331 4936 63340 4976
rect 63380 4936 63389 4976
rect 63331 4935 63389 4936
rect 64195 4976 64253 4977
rect 64195 4936 64204 4976
rect 64244 4936 64253 4976
rect 64195 4935 64253 4936
rect 65547 4976 65589 4985
rect 65547 4936 65548 4976
rect 65588 4936 65589 4976
rect 65547 4927 65589 4936
rect 65739 4976 65781 4985
rect 65739 4936 65740 4976
rect 65780 4936 65781 4976
rect 65739 4927 65781 4936
rect 65827 4976 65885 4977
rect 65827 4936 65836 4976
rect 65876 4936 65885 4976
rect 65827 4935 65885 4936
rect 66115 4976 66173 4977
rect 66115 4936 66124 4976
rect 66164 4936 66173 4976
rect 66115 4935 66173 4936
rect 66315 4976 66357 4985
rect 66315 4936 66316 4976
rect 66356 4936 66357 4976
rect 66315 4927 66357 4936
rect 66499 4976 66557 4977
rect 66499 4936 66508 4976
rect 66548 4936 66557 4976
rect 66499 4935 66557 4936
rect 66699 4976 66741 4985
rect 66699 4936 66700 4976
rect 66740 4936 66741 4976
rect 66699 4927 66741 4936
rect 68811 4976 68853 4985
rect 68811 4936 68812 4976
rect 68852 4936 68853 4976
rect 68811 4927 68853 4936
rect 69003 4976 69045 4985
rect 69003 4936 69004 4976
rect 69044 4936 69045 4976
rect 69003 4927 69045 4936
rect 69091 4976 69149 4977
rect 69091 4936 69100 4976
rect 69140 4936 69149 4976
rect 69091 4935 69149 4936
rect 71211 4976 71253 4985
rect 71211 4936 71212 4976
rect 71252 4936 71253 4976
rect 71211 4927 71253 4936
rect 71395 4976 71453 4977
rect 71395 4936 71404 4976
rect 71444 4936 71453 4976
rect 71395 4935 71453 4936
rect 71595 4976 71637 4985
rect 71595 4936 71596 4976
rect 71636 4936 71637 4976
rect 71595 4927 71637 4936
rect 71787 4976 71829 4985
rect 71787 4936 71788 4976
rect 71828 4936 71829 4976
rect 71787 4927 71829 4936
rect 71875 4976 71933 4977
rect 71875 4936 71884 4976
rect 71924 4936 71933 4976
rect 71875 4935 71933 4936
rect 75907 4976 75965 4977
rect 75907 4936 75916 4976
rect 75956 4936 75965 4976
rect 75907 4935 75965 4936
rect 76011 4976 76053 4985
rect 76011 4936 76012 4976
rect 76052 4936 76053 4976
rect 76011 4927 76053 4936
rect 76203 4976 76245 4985
rect 76203 4936 76204 4976
rect 76244 4936 76245 4976
rect 76203 4927 76245 4936
rect 76395 4976 76437 4985
rect 76395 4936 76396 4976
rect 76436 4936 76437 4976
rect 76395 4927 76437 4936
rect 76587 4976 76629 4985
rect 76587 4936 76588 4976
rect 76628 4936 76629 4976
rect 76587 4927 76629 4936
rect 76675 4976 76733 4977
rect 76675 4936 76684 4976
rect 76724 4936 76733 4976
rect 76675 4935 76733 4936
rect 77163 4976 77205 4985
rect 77163 4936 77164 4976
rect 77204 4936 77205 4976
rect 77163 4927 77205 4936
rect 77355 4976 77397 4985
rect 77355 4936 77356 4976
rect 77396 4936 77397 4976
rect 77355 4927 77397 4936
rect 77443 4976 77501 4977
rect 77443 4936 77452 4976
rect 77492 4936 77501 4976
rect 77443 4935 77501 4936
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 1411 4892 1469 4893
rect 1411 4852 1420 4892
rect 1460 4852 1469 4892
rect 1411 4851 1469 4852
rect 5547 4808 5589 4817
rect 5547 4768 5548 4808
rect 5588 4768 5589 4808
rect 5547 4759 5589 4768
rect 5931 4808 5973 4817
rect 5931 4768 5932 4808
rect 5972 4768 5973 4808
rect 5931 4759 5973 4768
rect 50091 4808 50133 4817
rect 50091 4768 50092 4808
rect 50132 4768 50133 4808
rect 50091 4759 50133 4768
rect 52875 4808 52917 4817
rect 52875 4768 52876 4808
rect 52916 4768 52917 4808
rect 52875 4759 52917 4768
rect 61515 4808 61557 4817
rect 61515 4768 61516 4808
rect 61556 4768 61557 4808
rect 61515 4759 61557 4768
rect 66891 4808 66933 4817
rect 66891 4768 66892 4808
rect 66932 4768 66933 4808
rect 66891 4759 66933 4768
rect 69483 4808 69525 4817
rect 69483 4768 69484 4808
rect 69524 4768 69525 4808
rect 69483 4759 69525 4768
rect 72363 4808 72405 4817
rect 72363 4768 72364 4808
rect 72404 4768 72405 4808
rect 72363 4759 72405 4768
rect 74475 4808 74517 4817
rect 74475 4768 74476 4808
rect 74516 4768 74517 4808
rect 74475 4759 74517 4768
rect 77835 4808 77877 4817
rect 77835 4768 77836 4808
rect 77876 4768 77877 4808
rect 77835 4759 77877 4768
rect 1227 4724 1269 4733
rect 1227 4684 1228 4724
rect 1268 4684 1269 4724
rect 1227 4675 1269 4684
rect 48067 4724 48125 4725
rect 48067 4684 48076 4724
rect 48116 4684 48125 4724
rect 48067 4683 48125 4684
rect 49131 4724 49173 4733
rect 49131 4684 49132 4724
rect 49172 4684 49173 4724
rect 49131 4675 49173 4684
rect 51531 4724 51573 4733
rect 51531 4684 51532 4724
rect 51572 4684 51573 4724
rect 51531 4675 51573 4684
rect 58531 4724 58589 4725
rect 58531 4684 58540 4724
rect 58580 4684 58589 4724
rect 58531 4683 58589 4684
rect 61219 4724 61277 4725
rect 61219 4684 61228 4724
rect 61268 4684 61277 4724
rect 61219 4683 61277 4684
rect 66219 4724 66261 4733
rect 66219 4684 66220 4724
rect 66260 4684 66261 4724
rect 66219 4675 66261 4684
rect 66603 4724 66645 4733
rect 66603 4684 66604 4724
rect 66644 4684 66645 4724
rect 66603 4675 66645 4684
rect 68811 4724 68853 4733
rect 68811 4684 68812 4724
rect 68852 4684 68853 4724
rect 68811 4675 68853 4684
rect 71307 4724 71349 4733
rect 71307 4684 71308 4724
rect 71348 4684 71349 4724
rect 71307 4675 71349 4684
rect 71595 4724 71637 4733
rect 71595 4684 71596 4724
rect 71636 4684 71637 4724
rect 71595 4675 71637 4684
rect 76395 4724 76437 4733
rect 76395 4684 76396 4724
rect 76436 4684 76437 4724
rect 76395 4675 76437 4684
rect 77163 4724 77205 4733
rect 77163 4684 77164 4724
rect 77204 4684 77205 4724
rect 77163 4675 77205 4684
rect 576 4556 79584 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 79584 4556
rect 576 4492 79584 4516
rect 2379 4388 2421 4397
rect 2379 4348 2380 4388
rect 2420 4348 2421 4388
rect 2379 4339 2421 4348
rect 52003 4388 52061 4389
rect 52003 4348 52012 4388
rect 52052 4348 52061 4388
rect 52003 4347 52061 4348
rect 66211 4388 66269 4389
rect 66211 4348 66220 4388
rect 66260 4348 66269 4388
rect 66211 4347 66269 4348
rect 651 4304 693 4313
rect 651 4264 652 4304
rect 692 4264 693 4304
rect 651 4255 693 4264
rect 1803 4304 1845 4313
rect 1803 4264 1804 4304
rect 1844 4264 1845 4304
rect 1803 4255 1845 4264
rect 4195 4304 4253 4305
rect 4195 4264 4204 4304
rect 4244 4264 4253 4304
rect 4195 4263 4253 4264
rect 5067 4304 5109 4313
rect 5067 4264 5068 4304
rect 5108 4264 5109 4304
rect 5067 4255 5109 4264
rect 7651 4304 7709 4305
rect 7651 4264 7660 4304
rect 7700 4264 7709 4304
rect 7651 4263 7709 4264
rect 54691 4304 54749 4305
rect 54691 4264 54700 4304
rect 54740 4264 54749 4304
rect 54691 4263 54749 4264
rect 55083 4304 55125 4313
rect 55083 4264 55084 4304
rect 55124 4264 55125 4304
rect 55083 4255 55125 4264
rect 56803 4304 56861 4305
rect 56803 4264 56812 4304
rect 56852 4264 56861 4304
rect 56803 4263 56861 4264
rect 57963 4304 58005 4313
rect 57963 4264 57964 4304
rect 58004 4264 58005 4304
rect 57963 4255 58005 4264
rect 60171 4304 60213 4313
rect 60171 4264 60172 4304
rect 60212 4264 60213 4304
rect 60171 4255 60213 4264
rect 68803 4304 68861 4305
rect 68803 4264 68812 4304
rect 68852 4264 68861 4304
rect 68803 4263 68861 4264
rect 74275 4304 74333 4305
rect 74275 4264 74284 4304
rect 74324 4264 74333 4304
rect 74275 4263 74333 4264
rect 76867 4304 76925 4305
rect 76867 4264 76876 4304
rect 76916 4264 76925 4304
rect 76867 4263 76925 4264
rect 79459 4304 79517 4305
rect 79459 4264 79468 4304
rect 79508 4264 79517 4304
rect 79459 4263 79517 4264
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 1219 4220 1277 4221
rect 1219 4180 1228 4220
rect 1268 4180 1277 4220
rect 1219 4179 1277 4180
rect 4491 4220 4533 4229
rect 4491 4180 4492 4220
rect 4532 4180 4533 4220
rect 4491 4171 4533 4180
rect 2379 4136 2421 4145
rect 2379 4096 2380 4136
rect 2420 4096 2421 4136
rect 2379 4087 2421 4096
rect 2571 4136 2613 4145
rect 2571 4096 2572 4136
rect 2612 4096 2613 4136
rect 2571 4087 2613 4096
rect 2659 4136 2717 4137
rect 2659 4096 2668 4136
rect 2708 4096 2717 4136
rect 3051 4136 3093 4145
rect 2659 4095 2717 4096
rect 2859 4094 2901 4103
rect 2859 4054 2860 4094
rect 2900 4054 2901 4094
rect 3051 4096 3052 4136
rect 3092 4096 3093 4136
rect 3051 4087 3093 4096
rect 3139 4136 3197 4137
rect 3139 4096 3148 4136
rect 3188 4096 3197 4136
rect 3139 4095 3197 4096
rect 3523 4136 3581 4137
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 3523 4095 3581 4096
rect 3819 4136 3861 4145
rect 3819 4096 3820 4136
rect 3860 4096 3861 4136
rect 3819 4087 3861 4096
rect 4395 4136 4437 4145
rect 4395 4096 4396 4136
rect 4436 4096 4437 4136
rect 4395 4087 4437 4096
rect 4579 4136 4637 4137
rect 4579 4096 4588 4136
rect 4628 4096 4637 4136
rect 4579 4095 4637 4096
rect 4771 4136 4829 4137
rect 4771 4096 4780 4136
rect 4820 4096 4829 4136
rect 4771 4095 4829 4096
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 5067 4136 5109 4145
rect 5067 4096 5068 4136
rect 5108 4096 5109 4136
rect 5067 4087 5109 4096
rect 5259 4136 5301 4145
rect 5259 4096 5260 4136
rect 5300 4096 5301 4136
rect 5259 4087 5301 4096
rect 5635 4136 5693 4137
rect 5635 4096 5644 4136
rect 5684 4096 5693 4136
rect 5635 4095 5693 4096
rect 6499 4136 6557 4137
rect 6499 4096 6508 4136
rect 6548 4096 6557 4136
rect 6499 4095 6557 4096
rect 47403 4136 47445 4145
rect 47403 4096 47404 4136
rect 47444 4096 47445 4136
rect 47403 4087 47445 4096
rect 47499 4136 47541 4145
rect 47499 4096 47500 4136
rect 47540 4096 47541 4136
rect 47499 4087 47541 4096
rect 47595 4136 47637 4145
rect 47595 4096 47596 4136
rect 47636 4096 47637 4136
rect 47595 4087 47637 4096
rect 47691 4136 47733 4145
rect 47691 4096 47692 4136
rect 47732 4096 47733 4136
rect 47691 4087 47733 4096
rect 49987 4136 50045 4137
rect 49987 4096 49996 4136
rect 50036 4096 50045 4136
rect 49987 4095 50045 4096
rect 50851 4136 50909 4137
rect 50851 4096 50860 4136
rect 50900 4096 50909 4136
rect 50851 4095 50909 4096
rect 52299 4136 52341 4145
rect 52299 4096 52300 4136
rect 52340 4096 52341 4136
rect 52299 4087 52341 4096
rect 52675 4136 52733 4137
rect 52675 4096 52684 4136
rect 52724 4096 52733 4136
rect 52675 4095 52733 4096
rect 53539 4136 53597 4137
rect 53539 4096 53548 4136
rect 53588 4096 53597 4136
rect 53539 4095 53597 4096
rect 55563 4136 55605 4145
rect 55563 4096 55564 4136
rect 55604 4096 55605 4136
rect 55563 4087 55605 4096
rect 55659 4136 55701 4145
rect 55659 4096 55660 4136
rect 55700 4096 55701 4136
rect 55659 4087 55701 4096
rect 55755 4136 55797 4145
rect 55755 4096 55756 4136
rect 55796 4096 55797 4136
rect 55755 4087 55797 4096
rect 55851 4136 55893 4145
rect 55851 4096 55852 4136
rect 55892 4096 55893 4136
rect 55851 4087 55893 4096
rect 56131 4136 56189 4137
rect 56131 4096 56140 4136
rect 56180 4096 56189 4136
rect 56131 4095 56189 4096
rect 56427 4136 56469 4145
rect 56427 4096 56428 4136
rect 56468 4096 56469 4136
rect 56427 4087 56469 4096
rect 57003 4136 57045 4145
rect 57003 4096 57004 4136
rect 57044 4096 57045 4136
rect 57003 4087 57045 4096
rect 57195 4136 57237 4145
rect 57195 4096 57196 4136
rect 57236 4096 57237 4136
rect 57195 4087 57237 4096
rect 57283 4136 57341 4137
rect 57283 4096 57292 4136
rect 57332 4096 57341 4136
rect 57283 4095 57341 4096
rect 57963 4136 58005 4145
rect 57963 4096 57964 4136
rect 58004 4096 58005 4136
rect 57963 4087 58005 4096
rect 58155 4136 58197 4145
rect 58155 4096 58156 4136
rect 58196 4096 58197 4136
rect 58155 4087 58197 4096
rect 58243 4136 58301 4137
rect 58243 4096 58252 4136
rect 58292 4096 58301 4136
rect 58243 4095 58301 4096
rect 58923 4136 58965 4145
rect 58923 4096 58924 4136
rect 58964 4096 58965 4136
rect 58923 4087 58965 4096
rect 59019 4136 59061 4145
rect 59019 4096 59020 4136
rect 59060 4096 59061 4136
rect 59019 4087 59061 4096
rect 59115 4136 59157 4145
rect 59115 4096 59116 4136
rect 59156 4096 59157 4136
rect 59115 4087 59157 4096
rect 59211 4136 59253 4145
rect 59211 4096 59212 4136
rect 59252 4096 59253 4136
rect 59211 4087 59253 4096
rect 63235 4136 63293 4137
rect 63235 4096 63244 4136
rect 63284 4096 63293 4136
rect 63235 4095 63293 4096
rect 64099 4136 64157 4137
rect 64099 4096 64108 4136
rect 64148 4096 64157 4136
rect 64099 4095 64157 4096
rect 65539 4136 65597 4137
rect 65539 4096 65548 4136
rect 65588 4096 65597 4136
rect 65539 4095 65597 4096
rect 65835 4136 65877 4145
rect 65835 4096 65836 4136
rect 65876 4096 65877 4136
rect 65835 4087 65877 4096
rect 66787 4136 66845 4137
rect 66787 4096 66796 4136
rect 66836 4096 66845 4136
rect 66787 4095 66845 4096
rect 67651 4136 67709 4137
rect 67651 4096 67660 4136
rect 67700 4096 67709 4136
rect 67651 4095 67709 4096
rect 69379 4136 69437 4137
rect 69379 4096 69388 4136
rect 69428 4096 69437 4136
rect 69379 4095 69437 4096
rect 70243 4136 70301 4137
rect 70243 4096 70252 4136
rect 70292 4096 70301 4136
rect 70243 4095 70301 4096
rect 71883 4136 71925 4145
rect 71883 4096 71884 4136
rect 71924 4096 71925 4136
rect 71883 4087 71925 4096
rect 72259 4136 72317 4137
rect 72259 4096 72268 4136
rect 72308 4096 72317 4136
rect 72259 4095 72317 4096
rect 73123 4136 73181 4137
rect 73123 4096 73132 4136
rect 73172 4096 73181 4136
rect 73123 4095 73181 4096
rect 74475 4136 74517 4145
rect 74475 4096 74476 4136
rect 74516 4096 74517 4136
rect 74475 4087 74517 4096
rect 74851 4136 74909 4137
rect 74851 4096 74860 4136
rect 74900 4096 74909 4136
rect 74851 4095 74909 4096
rect 75715 4136 75773 4137
rect 75715 4096 75724 4136
rect 75764 4096 75773 4136
rect 75715 4095 75773 4096
rect 77067 4136 77109 4145
rect 77067 4096 77068 4136
rect 77108 4096 77109 4136
rect 77067 4087 77109 4096
rect 77443 4136 77501 4137
rect 77443 4096 77452 4136
rect 77492 4096 77501 4136
rect 77443 4095 77501 4096
rect 78307 4136 78365 4137
rect 78307 4096 78316 4136
rect 78356 4096 78365 4136
rect 78307 4095 78365 4096
rect 2859 4045 2901 4054
rect 3915 4052 3957 4061
rect 3915 4012 3916 4052
rect 3956 4012 3957 4052
rect 3915 4003 3957 4012
rect 49611 4052 49653 4061
rect 49611 4012 49612 4052
rect 49652 4012 49653 4052
rect 49611 4003 49653 4012
rect 56523 4052 56565 4061
rect 56523 4012 56524 4052
rect 56564 4012 56565 4052
rect 56523 4003 56565 4012
rect 62859 4052 62901 4061
rect 62859 4012 62860 4052
rect 62900 4012 62901 4052
rect 62859 4003 62901 4012
rect 65931 4052 65973 4061
rect 65931 4012 65932 4052
rect 65972 4012 65973 4052
rect 65931 4003 65973 4012
rect 66411 4052 66453 4061
rect 66411 4012 66412 4052
rect 66452 4012 66453 4052
rect 66411 4003 66453 4012
rect 69003 4052 69045 4061
rect 69003 4012 69004 4052
rect 69044 4012 69045 4052
rect 69003 4003 69045 4012
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 2947 3968 3005 3969
rect 2947 3928 2956 3968
rect 2996 3928 3005 3968
rect 2947 3927 3005 3928
rect 52003 3968 52061 3969
rect 52003 3928 52012 3968
rect 52052 3928 52061 3968
rect 52003 3927 52061 3928
rect 57091 3968 57149 3969
rect 57091 3928 57100 3968
rect 57140 3928 57149 3968
rect 57091 3927 57149 3928
rect 65251 3968 65309 3969
rect 65251 3928 65260 3968
rect 65300 3928 65309 3968
rect 65251 3927 65309 3928
rect 71395 3968 71453 3969
rect 71395 3928 71404 3968
rect 71444 3928 71453 3968
rect 71395 3927 71453 3928
rect 576 3800 79584 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 79584 3800
rect 576 3736 79584 3760
rect 3715 3632 3773 3633
rect 3715 3592 3724 3632
rect 3764 3592 3773 3632
rect 3715 3591 3773 3592
rect 50179 3632 50237 3633
rect 50179 3592 50188 3632
rect 50228 3592 50237 3632
rect 50179 3591 50237 3592
rect 62083 3632 62141 3633
rect 62083 3592 62092 3632
rect 62132 3592 62141 3632
rect 62083 3591 62141 3592
rect 64003 3632 64061 3633
rect 64003 3592 64012 3632
rect 64052 3592 64061 3632
rect 64003 3591 64061 3592
rect 66211 3632 66269 3633
rect 66211 3592 66220 3632
rect 66260 3592 66269 3632
rect 66211 3591 66269 3592
rect 69283 3632 69341 3633
rect 69283 3592 69292 3632
rect 69332 3592 69341 3632
rect 69283 3591 69341 3592
rect 76099 3632 76157 3633
rect 76099 3592 76108 3632
rect 76148 3592 76157 3632
rect 76099 3591 76157 3592
rect 1323 3548 1365 3557
rect 1323 3508 1324 3548
rect 1364 3508 1365 3548
rect 1323 3499 1365 3508
rect 4395 3548 4437 3557
rect 4395 3508 4396 3548
rect 4436 3508 4437 3548
rect 4395 3499 4437 3508
rect 52011 3548 52053 3557
rect 52011 3508 52012 3548
rect 52052 3508 52053 3548
rect 52011 3499 52053 3508
rect 56139 3548 56181 3557
rect 56139 3508 56140 3548
rect 56180 3508 56181 3548
rect 56139 3499 56181 3508
rect 56715 3548 56757 3557
rect 56715 3508 56716 3548
rect 56756 3508 56757 3548
rect 56715 3499 56757 3508
rect 71403 3548 71445 3557
rect 71403 3508 71404 3548
rect 71444 3508 71445 3548
rect 71403 3499 71445 3508
rect 72171 3548 72213 3557
rect 72171 3508 72172 3548
rect 72212 3508 72213 3548
rect 72171 3499 72213 3508
rect 76779 3548 76821 3557
rect 76779 3508 76780 3548
rect 76820 3508 76821 3548
rect 76779 3499 76821 3508
rect 77355 3548 77397 3557
rect 77355 3508 77356 3548
rect 77396 3508 77397 3548
rect 77355 3499 77397 3508
rect 77739 3548 77781 3557
rect 77739 3508 77740 3548
rect 77780 3508 77781 3548
rect 77739 3499 77781 3508
rect 1699 3464 1757 3465
rect 1699 3424 1708 3464
rect 1748 3424 1757 3464
rect 1699 3423 1757 3424
rect 2563 3464 2621 3465
rect 2563 3424 2572 3464
rect 2612 3424 2621 3464
rect 2563 3423 2621 3424
rect 4299 3464 4341 3473
rect 4299 3424 4300 3464
rect 4340 3424 4341 3464
rect 4299 3415 4341 3424
rect 4483 3464 4541 3465
rect 4483 3424 4492 3464
rect 4532 3424 4541 3464
rect 4483 3423 4541 3424
rect 49987 3464 50045 3465
rect 49987 3424 49996 3464
rect 50036 3424 50045 3464
rect 49987 3423 50045 3424
rect 50091 3464 50133 3473
rect 50091 3424 50092 3464
rect 50132 3424 50133 3464
rect 50091 3415 50133 3424
rect 50283 3464 50325 3473
rect 50283 3424 50284 3464
rect 50324 3424 50325 3464
rect 50283 3415 50325 3424
rect 50571 3464 50613 3473
rect 50571 3424 50572 3464
rect 50612 3424 50613 3464
rect 50571 3415 50613 3424
rect 50667 3464 50709 3473
rect 50667 3424 50668 3464
rect 50708 3424 50709 3464
rect 50667 3415 50709 3424
rect 50763 3464 50805 3473
rect 50763 3424 50764 3464
rect 50804 3424 50805 3464
rect 50763 3415 50805 3424
rect 50859 3464 50901 3473
rect 50859 3424 50860 3464
rect 50900 3424 50901 3464
rect 50859 3415 50901 3424
rect 51619 3464 51677 3465
rect 51619 3424 51628 3464
rect 51668 3424 51677 3464
rect 51619 3423 51677 3424
rect 51915 3464 51957 3473
rect 51915 3424 51916 3464
rect 51956 3424 51957 3464
rect 51915 3415 51957 3424
rect 52491 3464 52533 3473
rect 52491 3424 52492 3464
rect 52532 3424 52533 3464
rect 52491 3415 52533 3424
rect 52675 3464 52733 3465
rect 52675 3424 52684 3464
rect 52724 3424 52733 3464
rect 52675 3423 52733 3424
rect 54883 3464 54941 3465
rect 54883 3424 54892 3464
rect 54932 3424 54941 3464
rect 54883 3423 54941 3424
rect 55747 3464 55805 3465
rect 55747 3424 55756 3464
rect 55796 3424 55805 3464
rect 55747 3423 55805 3424
rect 56611 3464 56669 3465
rect 56611 3424 56620 3464
rect 56660 3424 56669 3464
rect 56611 3423 56669 3424
rect 56811 3464 56853 3473
rect 56811 3424 56812 3464
rect 56852 3424 56853 3464
rect 56811 3415 56853 3424
rect 59299 3464 59357 3465
rect 59299 3424 59308 3464
rect 59348 3424 59357 3464
rect 59299 3423 59357 3424
rect 59499 3464 59541 3473
rect 59499 3424 59500 3464
rect 59540 3424 59541 3464
rect 59499 3415 59541 3424
rect 59691 3464 59733 3473
rect 59691 3424 59692 3464
rect 59732 3424 59733 3464
rect 59691 3415 59733 3424
rect 60067 3464 60125 3465
rect 60067 3424 60076 3464
rect 60116 3424 60125 3464
rect 60067 3423 60125 3424
rect 60931 3464 60989 3465
rect 60931 3424 60940 3464
rect 60980 3424 60989 3464
rect 60931 3423 60989 3424
rect 63811 3464 63869 3465
rect 63811 3424 63820 3464
rect 63860 3424 63869 3464
rect 63811 3423 63869 3424
rect 63915 3464 63957 3473
rect 63915 3424 63916 3464
rect 63956 3424 63957 3464
rect 63915 3415 63957 3424
rect 64107 3464 64149 3473
rect 64107 3424 64108 3464
rect 64148 3424 64149 3464
rect 64107 3415 64149 3424
rect 64299 3464 64341 3473
rect 64299 3424 64300 3464
rect 64340 3424 64341 3464
rect 64299 3415 64341 3424
rect 64395 3464 64437 3473
rect 64395 3424 64396 3464
rect 64436 3424 64437 3464
rect 64395 3415 64437 3424
rect 64491 3464 64533 3473
rect 64491 3424 64492 3464
rect 64532 3424 64533 3464
rect 64491 3415 64533 3424
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 66123 3464 66165 3473
rect 66123 3424 66124 3464
rect 66164 3424 66165 3464
rect 66123 3415 66165 3424
rect 66315 3464 66357 3473
rect 66315 3424 66316 3464
rect 66356 3424 66357 3464
rect 66315 3415 66357 3424
rect 66403 3464 66461 3465
rect 66403 3424 66412 3464
rect 66452 3424 66461 3464
rect 66403 3423 66461 3424
rect 68611 3464 68669 3465
rect 68611 3424 68620 3464
rect 68660 3424 68669 3464
rect 68611 3423 68669 3424
rect 68715 3464 68757 3473
rect 68715 3424 68716 3464
rect 68756 3424 68757 3464
rect 68715 3415 68757 3424
rect 68907 3464 68949 3473
rect 68907 3424 68908 3464
rect 68948 3424 68949 3464
rect 68907 3415 68949 3424
rect 69091 3464 69149 3465
rect 69091 3424 69100 3464
rect 69140 3424 69149 3464
rect 69091 3423 69149 3424
rect 69195 3464 69237 3473
rect 69195 3424 69196 3464
rect 69236 3424 69237 3464
rect 69195 3415 69237 3424
rect 69387 3464 69429 3473
rect 69387 3424 69388 3464
rect 69428 3424 69429 3464
rect 69387 3415 69429 3424
rect 69675 3464 69717 3473
rect 69675 3424 69676 3464
rect 69716 3424 69717 3464
rect 69675 3415 69717 3424
rect 69771 3464 69813 3473
rect 69771 3424 69772 3464
rect 69812 3424 69813 3464
rect 69771 3415 69813 3424
rect 69867 3464 69909 3473
rect 69867 3424 69868 3464
rect 69908 3424 69909 3464
rect 69867 3415 69909 3424
rect 69963 3464 70005 3473
rect 69963 3424 69964 3464
rect 70004 3424 70005 3464
rect 69963 3415 70005 3424
rect 70627 3464 70685 3465
rect 70627 3424 70636 3464
rect 70676 3424 70685 3464
rect 70627 3423 70685 3424
rect 70731 3464 70773 3473
rect 70731 3424 70732 3464
rect 70772 3424 70773 3464
rect 70731 3415 70773 3424
rect 70923 3464 70965 3473
rect 70923 3424 70924 3464
rect 70964 3424 70965 3464
rect 70923 3415 70965 3424
rect 71499 3464 71541 3473
rect 71499 3424 71500 3464
rect 71540 3424 71541 3464
rect 71499 3415 71541 3424
rect 71779 3464 71837 3465
rect 71779 3424 71788 3464
rect 71828 3424 71837 3464
rect 71779 3423 71837 3424
rect 72067 3464 72125 3465
rect 72067 3424 72076 3464
rect 72116 3424 72125 3464
rect 72067 3423 72125 3424
rect 72267 3464 72309 3473
rect 72267 3424 72268 3464
rect 72308 3424 72309 3464
rect 72267 3415 72309 3424
rect 72451 3464 72509 3465
rect 72451 3424 72460 3464
rect 72500 3424 72509 3464
rect 72451 3423 72509 3424
rect 72835 3464 72893 3465
rect 72835 3424 72844 3464
rect 72884 3424 72893 3464
rect 72835 3423 72893 3424
rect 73035 3464 73077 3473
rect 73035 3424 73036 3464
rect 73076 3424 73077 3464
rect 73035 3415 73077 3424
rect 75819 3464 75861 3473
rect 75819 3424 75820 3464
rect 75860 3424 75861 3464
rect 75819 3415 75861 3424
rect 75915 3464 75957 3473
rect 75915 3424 75916 3464
rect 75956 3424 75957 3464
rect 75915 3415 75957 3424
rect 76011 3464 76053 3473
rect 76011 3424 76012 3464
rect 76052 3424 76053 3464
rect 76011 3415 76053 3424
rect 76387 3464 76445 3465
rect 76387 3424 76396 3464
rect 76436 3424 76445 3464
rect 76387 3423 76445 3424
rect 76683 3464 76725 3473
rect 76683 3424 76684 3464
rect 76724 3424 76725 3464
rect 76683 3415 76725 3424
rect 77259 3464 77301 3473
rect 77259 3424 77260 3464
rect 77300 3424 77301 3464
rect 77259 3415 77301 3424
rect 77443 3464 77501 3465
rect 77443 3424 77452 3464
rect 77492 3424 77501 3464
rect 77443 3423 77501 3424
rect 77635 3464 77693 3465
rect 77635 3424 77644 3464
rect 77684 3424 77693 3464
rect 77635 3423 77693 3424
rect 77835 3464 77877 3473
rect 77835 3424 77836 3464
rect 77876 3424 77877 3464
rect 77835 3415 77877 3424
rect 1123 3380 1181 3381
rect 1123 3340 1132 3380
rect 1172 3340 1181 3380
rect 1123 3339 1181 3340
rect 63339 3338 63381 3347
rect 52291 3296 52349 3297
rect 52291 3256 52300 3296
rect 52340 3256 52349 3296
rect 52291 3255 52349 3256
rect 52587 3296 52629 3305
rect 52587 3256 52588 3296
rect 52628 3256 52629 3296
rect 63339 3298 63340 3338
rect 63380 3298 63381 3338
rect 63339 3289 63381 3298
rect 68907 3296 68949 3305
rect 52587 3247 52629 3256
rect 68907 3256 68908 3296
rect 68948 3256 68949 3296
rect 68907 3247 68949 3256
rect 71107 3296 71165 3297
rect 71107 3256 71116 3296
rect 71156 3256 71165 3296
rect 71107 3255 71165 3256
rect 77059 3296 77117 3297
rect 77059 3256 77068 3296
rect 77108 3256 77117 3296
rect 77059 3255 77117 3256
rect 939 3212 981 3221
rect 939 3172 940 3212
rect 980 3172 981 3212
rect 939 3163 981 3172
rect 53731 3212 53789 3213
rect 53731 3172 53740 3212
rect 53780 3172 53789 3212
rect 53731 3171 53789 3172
rect 59403 3212 59445 3221
rect 59403 3172 59404 3212
rect 59444 3172 59445 3212
rect 59403 3163 59445 3172
rect 70923 3212 70965 3221
rect 70923 3172 70924 3212
rect 70964 3172 70965 3212
rect 70923 3163 70965 3172
rect 72939 3212 72981 3221
rect 72939 3172 72940 3212
rect 72980 3172 72981 3212
rect 72939 3163 72981 3172
rect 576 3044 79584 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 79584 3044
rect 576 2980 79584 3004
rect 651 2876 693 2885
rect 651 2836 652 2876
rect 692 2836 693 2876
rect 651 2827 693 2836
rect 3051 2876 3093 2885
rect 3051 2836 3052 2876
rect 3092 2836 3093 2876
rect 3051 2827 3093 2836
rect 58827 2876 58869 2885
rect 58827 2836 58828 2876
rect 58868 2836 58869 2876
rect 58827 2827 58869 2836
rect 64011 2876 64053 2885
rect 64011 2836 64012 2876
rect 64052 2836 64053 2876
rect 64011 2827 64053 2836
rect 72651 2876 72693 2885
rect 72651 2836 72652 2876
rect 72692 2836 72693 2876
rect 72651 2827 72693 2836
rect 73315 2876 73373 2877
rect 73315 2836 73324 2876
rect 73364 2836 73373 2876
rect 73315 2835 73373 2836
rect 76203 2876 76245 2885
rect 76203 2836 76204 2876
rect 76244 2836 76245 2876
rect 76203 2827 76245 2836
rect 1515 2792 1557 2801
rect 1515 2752 1516 2792
rect 1556 2752 1557 2792
rect 1515 2743 1557 2752
rect 53931 2792 53973 2801
rect 53931 2752 53932 2792
rect 53972 2752 53973 2792
rect 53931 2743 53973 2752
rect 56907 2792 56949 2801
rect 56907 2752 56908 2792
rect 56948 2752 56949 2792
rect 56907 2743 56949 2752
rect 60067 2792 60125 2793
rect 60067 2752 60076 2792
rect 60116 2752 60125 2792
rect 60067 2751 60125 2752
rect 62187 2792 62229 2801
rect 62187 2752 62188 2792
rect 62228 2752 62229 2792
rect 62187 2743 62229 2752
rect 66507 2792 66549 2801
rect 66507 2752 66508 2792
rect 66548 2752 66549 2792
rect 66507 2743 66549 2752
rect 68715 2792 68757 2801
rect 68715 2752 68716 2792
rect 68756 2752 68757 2792
rect 68715 2743 68757 2752
rect 70923 2792 70965 2801
rect 70923 2752 70924 2792
rect 70964 2752 70965 2792
rect 70923 2743 70965 2752
rect 74667 2792 74709 2801
rect 74667 2752 74668 2792
rect 74708 2752 74709 2792
rect 74667 2743 74709 2752
rect 76011 2792 76053 2801
rect 76011 2752 76012 2792
rect 76052 2752 76053 2792
rect 76011 2743 76053 2752
rect 77443 2792 77501 2793
rect 77443 2752 77452 2792
rect 77492 2752 77501 2792
rect 77443 2751 77501 2752
rect 78219 2792 78261 2801
rect 78219 2752 78220 2792
rect 78260 2752 78261 2792
rect 78219 2743 78261 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 1219 2708 1277 2709
rect 1219 2668 1228 2708
rect 1268 2668 1277 2708
rect 1219 2667 1277 2668
rect 1699 2708 1757 2709
rect 1699 2668 1708 2708
rect 1748 2668 1757 2708
rect 1699 2667 1757 2668
rect 60363 2708 60405 2717
rect 60363 2668 60364 2708
rect 60404 2668 60405 2708
rect 60363 2659 60405 2668
rect 64779 2708 64821 2717
rect 64779 2668 64780 2708
rect 64820 2668 64821 2708
rect 64779 2659 64821 2668
rect 71691 2661 71733 2670
rect 2475 2624 2517 2633
rect 2475 2584 2476 2624
rect 2516 2584 2517 2624
rect 2475 2575 2517 2584
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2667 2624 2709 2633
rect 2667 2584 2668 2624
rect 2708 2584 2709 2624
rect 2667 2575 2709 2584
rect 2763 2624 2805 2633
rect 2763 2584 2764 2624
rect 2804 2584 2805 2624
rect 2763 2575 2805 2584
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 3051 2575 3093 2584
rect 3243 2624 3285 2633
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 3331 2624 3389 2625
rect 3331 2584 3340 2624
rect 3380 2584 3389 2624
rect 3331 2583 3389 2584
rect 55747 2624 55805 2625
rect 55747 2584 55756 2624
rect 55796 2584 55805 2624
rect 55747 2583 55805 2584
rect 55851 2624 55893 2633
rect 55851 2584 55852 2624
rect 55892 2584 55893 2624
rect 56331 2624 56373 2633
rect 55851 2575 55893 2584
rect 56043 2582 56085 2591
rect 56043 2542 56044 2582
rect 56084 2542 56085 2582
rect 56331 2584 56332 2624
rect 56372 2584 56373 2624
rect 56331 2575 56373 2584
rect 56523 2624 56565 2633
rect 56523 2584 56524 2624
rect 56564 2584 56565 2624
rect 56523 2575 56565 2584
rect 56611 2624 56669 2625
rect 56611 2584 56620 2624
rect 56660 2584 56669 2624
rect 56611 2583 56669 2584
rect 56803 2624 56861 2625
rect 56803 2584 56812 2624
rect 56852 2584 56861 2624
rect 56803 2583 56861 2584
rect 57003 2624 57045 2633
rect 57003 2584 57004 2624
rect 57044 2584 57045 2624
rect 57003 2575 57045 2584
rect 57187 2624 57245 2625
rect 57187 2584 57196 2624
rect 57236 2584 57245 2624
rect 57187 2583 57245 2584
rect 57291 2624 57333 2633
rect 57291 2584 57292 2624
rect 57332 2584 57333 2624
rect 57291 2575 57333 2584
rect 57483 2624 57525 2633
rect 57483 2584 57484 2624
rect 57524 2584 57525 2624
rect 57483 2575 57525 2584
rect 58827 2624 58869 2633
rect 58827 2584 58828 2624
rect 58868 2584 58869 2624
rect 58827 2575 58869 2584
rect 59019 2624 59061 2633
rect 59019 2584 59020 2624
rect 59060 2584 59061 2624
rect 59019 2575 59061 2584
rect 59107 2624 59165 2625
rect 59107 2584 59116 2624
rect 59156 2584 59165 2624
rect 59107 2583 59165 2584
rect 59395 2624 59453 2625
rect 59395 2584 59404 2624
rect 59444 2584 59453 2624
rect 59395 2583 59453 2584
rect 59691 2624 59733 2633
rect 59691 2584 59692 2624
rect 59732 2584 59733 2624
rect 59691 2575 59733 2584
rect 60267 2624 60309 2633
rect 60267 2584 60268 2624
rect 60308 2584 60309 2624
rect 60267 2575 60309 2584
rect 60451 2624 60509 2625
rect 60451 2584 60460 2624
rect 60500 2584 60509 2624
rect 60451 2583 60509 2584
rect 63715 2624 63773 2625
rect 63715 2584 63724 2624
rect 63764 2584 63773 2624
rect 63715 2583 63773 2584
rect 63819 2624 63861 2633
rect 63819 2584 63820 2624
rect 63860 2584 63861 2624
rect 63819 2575 63861 2584
rect 64011 2624 64053 2633
rect 64011 2584 64012 2624
rect 64052 2584 64053 2624
rect 64011 2575 64053 2584
rect 64203 2624 64245 2633
rect 64203 2584 64204 2624
rect 64244 2584 64245 2624
rect 64203 2575 64245 2584
rect 64395 2624 64437 2633
rect 64395 2584 64396 2624
rect 64436 2584 64437 2624
rect 64395 2575 64437 2584
rect 64483 2624 64541 2625
rect 64483 2584 64492 2624
rect 64532 2584 64541 2624
rect 64483 2583 64541 2584
rect 64675 2624 64733 2625
rect 64675 2584 64684 2624
rect 64724 2584 64733 2624
rect 64675 2583 64733 2584
rect 64875 2624 64917 2633
rect 64875 2584 64876 2624
rect 64916 2584 64917 2624
rect 64875 2575 64917 2584
rect 68235 2624 68277 2633
rect 68235 2584 68236 2624
rect 68276 2584 68277 2624
rect 68235 2575 68277 2584
rect 68331 2624 68373 2633
rect 68331 2584 68332 2624
rect 68372 2584 68373 2624
rect 68331 2575 68373 2584
rect 68427 2624 68469 2633
rect 68427 2584 68428 2624
rect 68468 2584 68469 2624
rect 68427 2575 68469 2584
rect 68619 2624 68661 2633
rect 68619 2584 68620 2624
rect 68660 2584 68661 2624
rect 68619 2575 68661 2584
rect 68803 2624 68861 2625
rect 68803 2584 68812 2624
rect 68852 2584 68861 2624
rect 68803 2583 68861 2584
rect 68995 2624 69053 2625
rect 68995 2584 69004 2624
rect 69044 2584 69053 2624
rect 68995 2583 69053 2584
rect 69195 2624 69237 2633
rect 69195 2584 69196 2624
rect 69236 2584 69237 2624
rect 69195 2575 69237 2584
rect 71107 2624 71165 2625
rect 71107 2584 71116 2624
rect 71156 2584 71165 2624
rect 71107 2583 71165 2584
rect 71211 2624 71253 2633
rect 71211 2584 71212 2624
rect 71252 2584 71253 2624
rect 71211 2575 71253 2584
rect 71403 2624 71445 2633
rect 71403 2584 71404 2624
rect 71444 2584 71445 2624
rect 71403 2575 71445 2584
rect 71595 2624 71637 2633
rect 71595 2584 71596 2624
rect 71636 2584 71637 2624
rect 71691 2621 71692 2661
rect 71732 2621 71733 2661
rect 71779 2666 71837 2667
rect 71779 2626 71788 2666
rect 71828 2626 71837 2666
rect 71779 2625 71837 2626
rect 71691 2612 71733 2621
rect 71883 2624 71925 2633
rect 71595 2575 71637 2584
rect 71883 2584 71884 2624
rect 71924 2584 71925 2624
rect 71883 2575 71925 2584
rect 72163 2624 72221 2625
rect 72163 2584 72172 2624
rect 72212 2584 72221 2624
rect 72163 2583 72221 2584
rect 73611 2624 73653 2633
rect 73611 2584 73612 2624
rect 73652 2584 73653 2624
rect 73611 2575 73653 2584
rect 73707 2624 73749 2633
rect 73707 2584 73708 2624
rect 73748 2584 73749 2624
rect 73707 2575 73749 2584
rect 73987 2624 74045 2625
rect 73987 2584 73996 2624
rect 74036 2584 74045 2624
rect 73987 2583 74045 2584
rect 74283 2624 74325 2633
rect 74283 2584 74284 2624
rect 74324 2584 74325 2624
rect 74283 2575 74325 2584
rect 74467 2624 74525 2625
rect 74467 2584 74476 2624
rect 74516 2584 74525 2624
rect 74467 2583 74525 2584
rect 76203 2624 76245 2633
rect 76203 2584 76204 2624
rect 76244 2584 76245 2624
rect 76203 2575 76245 2584
rect 76395 2624 76437 2633
rect 76395 2584 76396 2624
rect 76436 2584 76437 2624
rect 76395 2575 76437 2584
rect 76483 2624 76541 2625
rect 76483 2584 76492 2624
rect 76532 2584 76541 2624
rect 76483 2583 76541 2584
rect 76771 2624 76829 2625
rect 76771 2584 76780 2624
rect 76820 2584 76829 2624
rect 76771 2583 76829 2584
rect 77067 2624 77109 2633
rect 77067 2584 77068 2624
rect 77108 2584 77109 2624
rect 77067 2575 77109 2584
rect 77643 2624 77685 2633
rect 77643 2584 77644 2624
rect 77684 2584 77685 2624
rect 77643 2575 77685 2584
rect 77827 2624 77885 2625
rect 77827 2584 77836 2624
rect 77876 2584 77885 2624
rect 77827 2583 77885 2584
rect 56043 2533 56085 2542
rect 59787 2540 59829 2549
rect 59787 2500 59788 2540
rect 59828 2500 59829 2540
rect 59787 2491 59829 2500
rect 69099 2540 69141 2549
rect 69099 2500 69100 2540
rect 69140 2500 69141 2540
rect 69099 2491 69141 2500
rect 74379 2540 74421 2549
rect 74379 2500 74380 2540
rect 74420 2500 74421 2540
rect 74379 2491 74421 2500
rect 77163 2540 77205 2549
rect 77163 2500 77164 2540
rect 77204 2500 77205 2540
rect 77163 2491 77205 2500
rect 77739 2540 77781 2549
rect 77739 2500 77740 2540
rect 77780 2500 77781 2540
rect 77739 2491 77781 2500
rect 1035 2456 1077 2465
rect 1035 2416 1036 2456
rect 1076 2416 1077 2456
rect 1035 2407 1077 2416
rect 55939 2456 55997 2457
rect 55939 2416 55948 2456
rect 55988 2416 55997 2456
rect 55939 2415 55997 2416
rect 56419 2456 56477 2457
rect 56419 2416 56428 2456
rect 56468 2416 56477 2456
rect 56419 2415 56477 2416
rect 57379 2456 57437 2457
rect 57379 2416 57388 2456
rect 57428 2416 57437 2456
rect 57379 2415 57437 2416
rect 64291 2456 64349 2457
rect 64291 2416 64300 2456
rect 64340 2416 64349 2456
rect 64291 2415 64349 2416
rect 68131 2456 68189 2457
rect 68131 2416 68140 2456
rect 68180 2416 68189 2456
rect 68131 2415 68189 2416
rect 71299 2456 71357 2457
rect 71299 2416 71308 2456
rect 71348 2416 71357 2456
rect 71299 2415 71357 2416
rect 72651 2456 72693 2465
rect 72651 2416 72652 2456
rect 72692 2416 72693 2456
rect 72651 2407 72693 2416
rect 576 2288 79584 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 79584 2288
rect 576 2224 79584 2248
rect 55843 2120 55901 2121
rect 55843 2080 55852 2120
rect 55892 2080 55901 2120
rect 55843 2079 55901 2080
rect 61603 2120 61661 2121
rect 61603 2080 61612 2120
rect 61652 2080 61661 2120
rect 61603 2079 61661 2080
rect 66883 2120 66941 2121
rect 66883 2080 66892 2120
rect 66932 2080 66941 2120
rect 66883 2079 66941 2080
rect 71203 2120 71261 2121
rect 71203 2080 71212 2120
rect 71252 2080 71261 2120
rect 71203 2079 71261 2080
rect 73795 2120 73853 2121
rect 73795 2080 73804 2120
rect 73844 2080 73853 2120
rect 73795 2079 73853 2080
rect 56619 2036 56661 2045
rect 56619 1996 56620 2036
rect 56660 1996 56661 2036
rect 56619 1987 56661 1996
rect 64491 2036 64533 2045
rect 64491 1996 64492 2036
rect 64532 1996 64533 2036
rect 64491 1987 64533 1996
rect 71403 2036 71445 2045
rect 71403 1996 71404 2036
rect 71444 1996 71445 2036
rect 71403 1987 71445 1996
rect 53451 1952 53493 1961
rect 53451 1912 53452 1952
rect 53492 1912 53493 1952
rect 53451 1903 53493 1912
rect 53827 1952 53885 1953
rect 53827 1912 53836 1952
rect 53876 1912 53885 1952
rect 53827 1911 53885 1912
rect 54691 1952 54749 1953
rect 54691 1912 54700 1952
rect 54740 1912 54749 1952
rect 54691 1911 54749 1912
rect 56043 1952 56085 1961
rect 56043 1912 56044 1952
rect 56084 1912 56085 1952
rect 56043 1903 56085 1912
rect 56235 1952 56277 1961
rect 56235 1912 56236 1952
rect 56276 1912 56277 1952
rect 56235 1903 56277 1912
rect 56323 1952 56381 1953
rect 56323 1912 56332 1952
rect 56372 1912 56381 1952
rect 56323 1911 56381 1912
rect 56995 1952 57053 1953
rect 56995 1912 57004 1952
rect 57044 1912 57053 1952
rect 56995 1911 57053 1912
rect 57859 1952 57917 1953
rect 57859 1912 57868 1952
rect 57908 1912 57917 1952
rect 57859 1911 57917 1912
rect 59211 1952 59253 1961
rect 59211 1912 59212 1952
rect 59252 1912 59253 1952
rect 59211 1903 59253 1912
rect 59587 1952 59645 1953
rect 59587 1912 59596 1952
rect 59636 1912 59645 1952
rect 59587 1911 59645 1912
rect 60451 1952 60509 1953
rect 60451 1912 60460 1952
rect 60500 1912 60509 1952
rect 60451 1911 60509 1912
rect 61803 1952 61845 1961
rect 61803 1912 61804 1952
rect 61844 1912 61845 1952
rect 61803 1903 61845 1912
rect 62179 1952 62237 1953
rect 62179 1912 62188 1952
rect 62228 1912 62237 1952
rect 62179 1911 62237 1912
rect 63043 1952 63101 1953
rect 63043 1912 63052 1952
rect 63092 1912 63101 1952
rect 63043 1911 63101 1912
rect 64867 1952 64925 1953
rect 64867 1912 64876 1952
rect 64916 1912 64925 1952
rect 64867 1911 64925 1912
rect 65731 1952 65789 1953
rect 65731 1912 65740 1952
rect 65780 1912 65789 1952
rect 65731 1911 65789 1912
rect 67371 1952 67413 1961
rect 67371 1912 67372 1952
rect 67412 1912 67413 1952
rect 67371 1903 67413 1912
rect 67563 1952 67605 1961
rect 67563 1912 67564 1952
rect 67604 1912 67605 1952
rect 67563 1903 67605 1912
rect 67651 1952 67709 1953
rect 67651 1912 67660 1952
rect 67700 1912 67709 1952
rect 67651 1911 67709 1912
rect 67939 1952 67997 1953
rect 67939 1912 67948 1952
rect 67988 1912 67997 1952
rect 67939 1911 67997 1912
rect 68235 1952 68277 1961
rect 68235 1912 68236 1952
rect 68276 1912 68277 1952
rect 68235 1903 68277 1912
rect 68331 1952 68373 1961
rect 68331 1912 68332 1952
rect 68372 1912 68373 1952
rect 68331 1903 68373 1912
rect 68811 1952 68853 1961
rect 68811 1912 68812 1952
rect 68852 1912 68853 1952
rect 68811 1903 68853 1912
rect 69187 1952 69245 1953
rect 69187 1912 69196 1952
rect 69236 1912 69245 1952
rect 69187 1911 69245 1912
rect 70051 1952 70109 1953
rect 70051 1912 70060 1952
rect 70100 1912 70109 1952
rect 70051 1911 70109 1912
rect 71779 1952 71837 1953
rect 71779 1912 71788 1952
rect 71828 1912 71837 1952
rect 71779 1911 71837 1912
rect 72643 1952 72701 1953
rect 72643 1912 72652 1952
rect 72692 1912 72701 1952
rect 72643 1911 72701 1912
rect 73995 1952 74037 1961
rect 73995 1912 73996 1952
rect 74036 1912 74037 1952
rect 73995 1903 74037 1912
rect 74187 1952 74229 1961
rect 74187 1912 74188 1952
rect 74228 1912 74229 1952
rect 74187 1903 74229 1912
rect 74275 1952 74333 1953
rect 74275 1912 74284 1952
rect 74324 1912 74333 1952
rect 74275 1911 74333 1912
rect 74563 1952 74621 1953
rect 74563 1912 74572 1952
rect 74612 1912 74621 1952
rect 74563 1911 74621 1912
rect 74667 1952 74709 1961
rect 74667 1912 74668 1952
rect 74708 1912 74709 1952
rect 74667 1903 74709 1912
rect 74859 1952 74901 1961
rect 74859 1912 74860 1952
rect 74900 1912 74901 1952
rect 74859 1903 74901 1912
rect 75139 1952 75197 1953
rect 75139 1912 75148 1952
rect 75188 1912 75197 1952
rect 75139 1911 75197 1912
rect 75243 1952 75285 1961
rect 75243 1912 75244 1952
rect 75284 1912 75285 1952
rect 75243 1903 75285 1912
rect 75435 1952 75477 1961
rect 75435 1912 75436 1952
rect 75476 1912 75477 1952
rect 75435 1903 75477 1912
rect 75627 1952 75669 1961
rect 75627 1912 75628 1952
rect 75668 1912 75669 1952
rect 75627 1903 75669 1912
rect 76003 1952 76061 1953
rect 76003 1912 76012 1952
rect 76052 1912 76061 1952
rect 76003 1911 76061 1912
rect 76867 1952 76925 1953
rect 76867 1912 76876 1952
rect 76916 1912 76925 1952
rect 76867 1911 76925 1912
rect 78219 1952 78261 1961
rect 78219 1912 78220 1952
rect 78260 1912 78261 1952
rect 78219 1903 78261 1912
rect 78411 1952 78453 1961
rect 78411 1912 78412 1952
rect 78452 1912 78453 1952
rect 78411 1903 78453 1912
rect 78499 1952 78557 1953
rect 78499 1912 78508 1952
rect 78548 1912 78557 1952
rect 78499 1911 78557 1912
rect 78691 1952 78749 1953
rect 78691 1912 78700 1952
rect 78740 1912 78749 1952
rect 78691 1911 78749 1912
rect 78891 1952 78933 1961
rect 78891 1912 78892 1952
rect 78932 1912 78933 1952
rect 78891 1903 78933 1912
rect 56043 1784 56085 1793
rect 56043 1744 56044 1784
rect 56084 1744 56085 1784
rect 56043 1735 56085 1744
rect 68611 1784 68669 1785
rect 68611 1744 68620 1784
rect 68660 1744 68669 1784
rect 68611 1743 68669 1744
rect 74859 1784 74901 1793
rect 74859 1744 74860 1784
rect 74900 1744 74901 1784
rect 74859 1735 74901 1744
rect 75435 1784 75477 1793
rect 75435 1744 75436 1784
rect 75476 1744 75477 1784
rect 75435 1735 75477 1744
rect 78795 1784 78837 1793
rect 78795 1744 78796 1784
rect 78836 1744 78837 1784
rect 78795 1735 78837 1744
rect 59011 1700 59069 1701
rect 59011 1660 59020 1700
rect 59060 1660 59069 1700
rect 59011 1659 59069 1660
rect 61603 1700 61661 1701
rect 61603 1660 61612 1700
rect 61652 1660 61661 1700
rect 61603 1659 61661 1660
rect 64195 1700 64253 1701
rect 64195 1660 64204 1700
rect 64244 1660 64253 1700
rect 64195 1659 64253 1660
rect 67371 1700 67413 1709
rect 67371 1660 67372 1700
rect 67412 1660 67413 1700
rect 67371 1651 67413 1660
rect 73995 1700 74037 1709
rect 73995 1660 73996 1700
rect 74036 1660 74037 1700
rect 73995 1651 74037 1660
rect 78019 1700 78077 1701
rect 78019 1660 78028 1700
rect 78068 1660 78077 1700
rect 78019 1659 78077 1660
rect 78219 1700 78261 1709
rect 78219 1660 78220 1700
rect 78260 1660 78261 1700
rect 78219 1651 78261 1660
rect 576 1532 79584 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 79584 1532
rect 576 1468 79584 1492
rect 56803 1364 56861 1365
rect 56803 1324 56812 1364
rect 56852 1324 56861 1364
rect 56803 1323 56861 1324
rect 58923 1364 58965 1373
rect 58923 1324 58924 1364
rect 58964 1324 58965 1364
rect 58923 1315 58965 1324
rect 62475 1364 62517 1373
rect 62475 1324 62476 1364
rect 62516 1324 62517 1364
rect 62475 1315 62517 1324
rect 68419 1364 68477 1365
rect 68419 1324 68428 1364
rect 68468 1324 68477 1364
rect 68419 1323 68477 1324
rect 68907 1364 68949 1373
rect 68907 1324 68908 1364
rect 68948 1324 68949 1364
rect 68907 1315 68949 1324
rect 70155 1364 70197 1373
rect 70155 1324 70156 1364
rect 70196 1324 70197 1364
rect 70155 1315 70197 1324
rect 71883 1364 71925 1373
rect 71883 1324 71884 1364
rect 71924 1324 71925 1364
rect 71883 1315 71925 1324
rect 75619 1364 75677 1365
rect 75619 1324 75628 1364
rect 75668 1324 75677 1364
rect 75619 1323 75677 1324
rect 77059 1364 77117 1365
rect 77059 1324 77068 1364
rect 77108 1324 77117 1364
rect 77059 1323 77117 1324
rect 57099 1280 57141 1289
rect 57099 1240 57100 1280
rect 57140 1240 57141 1280
rect 57099 1231 57141 1240
rect 57387 1280 57429 1289
rect 57387 1240 57388 1280
rect 57428 1240 57429 1280
rect 57387 1231 57429 1240
rect 60843 1280 60885 1289
rect 60843 1240 60844 1280
rect 60884 1240 60885 1280
rect 60843 1231 60885 1240
rect 61995 1280 62037 1289
rect 61995 1240 61996 1280
rect 62036 1240 62037 1280
rect 61995 1231 62037 1240
rect 64483 1280 64541 1281
rect 64483 1240 64492 1280
rect 64532 1240 64541 1280
rect 64483 1239 64541 1240
rect 64779 1280 64821 1289
rect 64779 1240 64780 1280
rect 64820 1240 64821 1280
rect 64779 1231 64821 1240
rect 65067 1280 65109 1289
rect 65067 1240 65068 1280
rect 65108 1240 65109 1280
rect 65067 1231 65109 1240
rect 69387 1280 69429 1289
rect 69387 1240 69388 1280
rect 69428 1240 69429 1280
rect 69387 1231 69429 1240
rect 55467 1112 55509 1121
rect 55467 1072 55468 1112
rect 55508 1072 55509 1112
rect 55467 1063 55509 1072
rect 55563 1112 55605 1121
rect 55563 1072 55564 1112
rect 55604 1072 55605 1112
rect 55563 1063 55605 1072
rect 55659 1112 55701 1121
rect 55659 1072 55660 1112
rect 55700 1072 55701 1112
rect 55659 1063 55701 1072
rect 55755 1112 55797 1121
rect 55755 1072 55756 1112
rect 55796 1072 55797 1112
rect 55755 1063 55797 1072
rect 56131 1112 56189 1113
rect 56131 1072 56140 1112
rect 56180 1072 56189 1112
rect 56131 1071 56189 1072
rect 56427 1112 56469 1121
rect 56427 1072 56428 1112
rect 56468 1072 56469 1112
rect 56427 1063 56469 1072
rect 56523 1112 56565 1121
rect 56523 1072 56524 1112
rect 56564 1072 56565 1112
rect 56523 1063 56565 1072
rect 56995 1112 57053 1113
rect 56995 1072 57004 1112
rect 57044 1072 57053 1112
rect 56995 1071 57053 1072
rect 57195 1112 57237 1121
rect 57195 1072 57196 1112
rect 57236 1072 57237 1112
rect 57195 1063 57237 1072
rect 58627 1112 58685 1113
rect 58627 1072 58636 1112
rect 58676 1072 58685 1112
rect 58627 1071 58685 1072
rect 58731 1112 58773 1121
rect 58731 1072 58732 1112
rect 58772 1072 58773 1112
rect 58731 1063 58773 1072
rect 58923 1112 58965 1121
rect 58923 1072 58924 1112
rect 58964 1072 58965 1112
rect 58923 1063 58965 1072
rect 59107 1112 59165 1113
rect 59107 1072 59116 1112
rect 59156 1072 59165 1112
rect 59107 1071 59165 1072
rect 60067 1112 60125 1113
rect 60067 1072 60076 1112
rect 60116 1072 60125 1112
rect 60067 1071 60125 1072
rect 60459 1112 60501 1121
rect 60459 1072 60460 1112
rect 60500 1072 60501 1112
rect 60459 1063 60501 1072
rect 60555 1112 60597 1121
rect 60555 1072 60556 1112
rect 60596 1072 60597 1112
rect 60555 1063 60597 1072
rect 60651 1112 60693 1121
rect 60651 1072 60652 1112
rect 60692 1072 60693 1112
rect 60651 1063 60693 1072
rect 61699 1112 61757 1113
rect 61699 1072 61708 1112
rect 61748 1072 61757 1112
rect 61699 1071 61757 1072
rect 61803 1112 61845 1121
rect 61803 1072 61804 1112
rect 61844 1072 61845 1112
rect 61803 1063 61845 1072
rect 61995 1112 62037 1121
rect 61995 1072 61996 1112
rect 62036 1072 62037 1112
rect 61995 1063 62037 1072
rect 62179 1112 62237 1113
rect 62179 1072 62188 1112
rect 62228 1072 62237 1112
rect 62179 1071 62237 1072
rect 62283 1112 62325 1121
rect 62283 1072 62284 1112
rect 62324 1072 62325 1112
rect 62283 1063 62325 1072
rect 62475 1112 62517 1121
rect 62475 1072 62476 1112
rect 62516 1072 62517 1112
rect 62475 1063 62517 1072
rect 62667 1112 62709 1121
rect 62667 1072 62668 1112
rect 62708 1072 62709 1112
rect 62667 1063 62709 1072
rect 62763 1112 62805 1121
rect 62763 1072 62764 1112
rect 62804 1072 62805 1112
rect 62763 1063 62805 1072
rect 62859 1112 62901 1121
rect 62859 1072 62860 1112
rect 62900 1072 62901 1112
rect 62859 1063 62901 1072
rect 62955 1112 62997 1121
rect 62955 1072 62956 1112
rect 62996 1072 62997 1112
rect 62955 1063 62997 1072
rect 63811 1112 63869 1113
rect 63811 1072 63820 1112
rect 63860 1072 63869 1112
rect 63811 1071 63869 1072
rect 64107 1112 64149 1121
rect 64107 1072 64108 1112
rect 64148 1072 64149 1112
rect 64107 1063 64149 1072
rect 64683 1112 64725 1121
rect 64683 1072 64684 1112
rect 64724 1072 64725 1112
rect 64683 1063 64725 1072
rect 64867 1112 64925 1113
rect 64867 1072 64876 1112
rect 64916 1072 64925 1112
rect 64867 1071 64925 1072
rect 66027 1112 66069 1121
rect 66027 1072 66028 1112
rect 66068 1072 66069 1112
rect 66027 1063 66069 1072
rect 66403 1112 66461 1113
rect 66403 1072 66412 1112
rect 66452 1072 66461 1112
rect 66403 1071 66461 1072
rect 67267 1112 67325 1113
rect 67267 1072 67276 1112
rect 67316 1072 67325 1112
rect 67267 1071 67325 1072
rect 68611 1112 68669 1113
rect 68611 1072 68620 1112
rect 68660 1072 68669 1112
rect 68611 1071 68669 1072
rect 68715 1112 68757 1121
rect 68715 1072 68716 1112
rect 68756 1072 68757 1112
rect 68715 1063 68757 1072
rect 68907 1112 68949 1121
rect 68907 1072 68908 1112
rect 68948 1072 68949 1112
rect 68907 1063 68949 1072
rect 70731 1112 70773 1121
rect 70731 1072 70732 1112
rect 70772 1072 70773 1112
rect 70731 1063 70773 1072
rect 71203 1112 71261 1113
rect 71203 1072 71212 1112
rect 71252 1072 71261 1112
rect 71203 1071 71261 1072
rect 72547 1112 72605 1113
rect 72547 1072 72556 1112
rect 72596 1072 72605 1112
rect 72547 1071 72605 1072
rect 73227 1112 73269 1121
rect 73227 1072 73228 1112
rect 73268 1072 73269 1112
rect 73227 1063 73269 1072
rect 73603 1112 73661 1113
rect 73603 1072 73612 1112
rect 73652 1072 73661 1112
rect 73603 1071 73661 1072
rect 74467 1112 74525 1113
rect 74467 1072 74476 1112
rect 74516 1072 74525 1112
rect 74467 1071 74525 1072
rect 76011 1112 76053 1121
rect 76011 1072 76012 1112
rect 76052 1072 76053 1112
rect 76011 1063 76053 1072
rect 76107 1112 76149 1121
rect 76107 1072 76108 1112
rect 76148 1072 76149 1112
rect 76107 1063 76149 1072
rect 76203 1112 76245 1121
rect 76203 1072 76204 1112
rect 76244 1072 76245 1112
rect 76203 1063 76245 1072
rect 78211 1112 78269 1113
rect 78211 1072 78220 1112
rect 78260 1072 78269 1112
rect 78211 1071 78269 1072
rect 79075 1112 79133 1113
rect 79075 1072 79084 1112
rect 79124 1072 79133 1112
rect 79075 1071 79133 1072
rect 79467 1112 79509 1121
rect 79467 1072 79468 1112
rect 79508 1072 79509 1112
rect 79467 1063 79509 1072
rect 64203 1028 64245 1037
rect 64203 988 64204 1028
rect 64244 988 64245 1028
rect 64203 979 64245 988
rect 60355 944 60413 945
rect 60355 904 60364 944
rect 60404 904 60413 944
rect 60355 903 60413 904
rect 75907 944 75965 945
rect 75907 904 75916 944
rect 75956 904 75965 944
rect 75907 903 75965 904
rect 576 776 79584 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 79584 776
rect 576 712 79584 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 64108 38284 64148 38324
rect 58060 38200 58100 38240
rect 58252 38200 58292 38240
rect 58348 38200 58388 38240
rect 59404 38200 59444 38240
rect 63532 38200 63572 38240
rect 63724 38200 63764 38240
rect 63820 38200 63860 38240
rect 64012 38200 64052 38240
rect 64204 38200 64244 38240
rect 67468 38200 67508 38240
rect 68044 38200 68084 38240
rect 68140 38200 68180 38240
rect 68236 38200 68276 38240
rect 68332 38200 68372 38240
rect 68716 38200 68756 38240
rect 68812 38200 68852 38240
rect 69004 38200 69044 38240
rect 70156 38200 70196 38240
rect 71404 38200 71444 38240
rect 72748 38200 72788 38240
rect 76876 38200 76916 38240
rect 77164 38200 77204 38240
rect 77260 38200 77300 38240
rect 652 38116 692 38156
rect 57292 38116 57332 38156
rect 57676 38116 57716 38156
rect 59980 38116 60020 38156
rect 67852 38116 67892 38156
rect 69388 38116 69428 38156
rect 70636 38116 70676 38156
rect 56428 38032 56468 38072
rect 57868 38032 57908 38072
rect 60172 38032 60212 38072
rect 61900 38032 61940 38072
rect 64588 38032 64628 38072
rect 66220 38032 66260 38072
rect 71980 38032 72020 38072
rect 73996 38032 74036 38072
rect 76012 38032 76052 38072
rect 844 37948 884 37988
rect 57484 37948 57524 37988
rect 58060 37948 58100 37988
rect 58828 37948 58868 37988
rect 59788 37948 59828 37988
rect 63532 37948 63572 37988
rect 67660 37948 67700 37988
rect 69004 37948 69044 37988
rect 73036 37948 73076 37988
rect 77548 37948 77588 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 67756 37612 67796 37652
rect 54892 37528 54932 37568
rect 78508 37528 78548 37568
rect 67564 37444 67604 37484
rect 55468 37360 55508 37400
rect 55660 37360 55700 37400
rect 55756 37360 55796 37400
rect 55948 37360 55988 37400
rect 56332 37360 56372 37400
rect 57196 37360 57236 37400
rect 58540 37360 58580 37400
rect 58636 37360 58676 37400
rect 58732 37360 58772 37400
rect 59500 37360 59540 37400
rect 60364 37360 60404 37400
rect 62092 37360 62132 37400
rect 62956 37360 62996 37400
rect 64300 37360 64340 37400
rect 64684 37360 64724 37400
rect 65548 37360 65588 37400
rect 67084 37360 67124 37400
rect 67276 37360 67316 37400
rect 67372 37360 67412 37400
rect 68044 37360 68084 37400
rect 68332 37360 68372 37400
rect 69100 37360 69140 37400
rect 69484 37360 69524 37400
rect 70348 37360 70388 37400
rect 72748 37360 72788 37400
rect 72844 37360 72884 37400
rect 72940 37360 72980 37400
rect 73228 37360 73268 37400
rect 73516 37360 73556 37400
rect 73708 37360 73748 37400
rect 59116 37276 59156 37316
rect 61708 37276 61748 37316
rect 68428 37276 68468 37316
rect 73036 37276 73076 37316
rect 73420 37318 73460 37358
rect 73900 37360 73940 37400
rect 73996 37360 74036 37400
rect 74284 37360 74324 37400
rect 74476 37360 74516 37400
rect 74572 37360 74612 37400
rect 75052 37360 75092 37400
rect 75148 37360 75188 37400
rect 75244 37360 75284 37400
rect 75916 37360 75956 37400
rect 76780 37360 76820 37400
rect 78124 37360 78164 37400
rect 78316 37360 78356 37400
rect 74380 37276 74420 37316
rect 75532 37276 75572 37316
rect 78220 37276 78260 37316
rect 55564 37192 55604 37232
rect 58348 37192 58388 37232
rect 58828 37192 58868 37232
rect 61516 37192 61556 37232
rect 64108 37192 64148 37232
rect 66700 37192 66740 37232
rect 67180 37192 67220 37232
rect 67756 37192 67796 37232
rect 71500 37192 71540 37232
rect 73324 37192 73364 37232
rect 73804 37192 73844 37232
rect 75340 37192 75380 37232
rect 77932 37192 77972 37232
rect 68716 37150 68756 37190
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 57100 36856 57140 36896
rect 59212 36856 59252 36896
rect 60268 36856 60308 36896
rect 61996 36856 62036 36896
rect 68140 36856 68180 36896
rect 76204 36856 76244 36896
rect 79468 36856 79508 36896
rect 54412 36772 54452 36812
rect 59692 36772 59732 36812
rect 63532 36772 63572 36812
rect 69004 36772 69044 36812
rect 69388 36772 69428 36812
rect 73324 36772 73364 36812
rect 73516 36772 73556 36812
rect 54796 36688 54836 36728
rect 55660 36688 55700 36728
rect 57004 36688 57044 36728
rect 57196 36688 57236 36728
rect 57292 36688 57332 36728
rect 58252 36688 58292 36728
rect 58540 36688 58580 36728
rect 58636 36688 58676 36728
rect 59116 36688 59156 36728
rect 59308 36688 59348 36728
rect 59404 36688 59444 36728
rect 59596 36688 59636 36728
rect 59788 36688 59828 36728
rect 60172 36688 60212 36728
rect 60364 36688 60404 36728
rect 60460 36688 60500 36728
rect 61420 36688 61460 36728
rect 61516 36688 61556 36728
rect 61612 36688 61652 36728
rect 61708 36688 61748 36728
rect 61900 36688 61940 36728
rect 62092 36688 62132 36728
rect 62188 36688 62228 36728
rect 63148 36688 63188 36728
rect 63436 36688 63476 36728
rect 64012 36688 64052 36728
rect 64204 36688 64244 36728
rect 65740 36688 65780 36728
rect 66124 36688 66164 36728
rect 66988 36688 67028 36728
rect 68428 36688 68468 36728
rect 68620 36688 68660 36728
rect 68716 36688 68756 36728
rect 68908 36688 68948 36728
rect 69095 36665 69135 36705
rect 69292 36688 69332 36728
rect 69484 36688 69524 36728
rect 72076 36688 72116 36728
rect 72940 36688 72980 36728
rect 73900 36688 73940 36728
rect 74764 36688 74804 36728
rect 76108 36688 76148 36728
rect 76300 36688 76340 36728
rect 76396 36688 76436 36728
rect 76588 36688 76628 36728
rect 76780 36688 76820 36728
rect 76876 36688 76916 36728
rect 77068 36688 77108 36728
rect 77452 36688 77492 36728
rect 78316 36688 78356 36728
rect 63820 36520 63860 36560
rect 64108 36520 64148 36560
rect 69676 36520 69716 36560
rect 76588 36520 76628 36560
rect 56812 36436 56852 36476
rect 58924 36436 58964 36476
rect 68428 36436 68468 36476
rect 70924 36436 70964 36476
rect 75916 36436 75956 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 73708 36100 73748 36140
rect 74092 36100 74132 36140
rect 76492 36100 76532 36140
rect 77548 36100 77588 36140
rect 49132 36016 49172 36056
rect 60268 36016 60308 36056
rect 69484 36016 69524 36056
rect 74668 36016 74708 36056
rect 50956 35932 50996 35972
rect 56812 35932 56852 35972
rect 73420 35974 73460 36014
rect 77836 36016 77876 36056
rect 58924 35932 58964 35972
rect 51244 35848 51284 35888
rect 51436 35848 51476 35888
rect 52396 35848 52436 35888
rect 53260 35837 53300 35877
rect 55756 35848 55796 35888
rect 55852 35848 55892 35888
rect 55948 35848 55988 35888
rect 56044 35848 56084 35888
rect 56236 35848 56276 35888
rect 56428 35848 56468 35888
rect 58828 35848 58868 35888
rect 59020 35848 59060 35888
rect 61324 35848 61364 35888
rect 61516 35848 61556 35888
rect 61612 35848 61652 35888
rect 61900 35848 61940 35888
rect 61996 35848 62036 35888
rect 62092 35848 62132 35888
rect 64588 35848 64628 35888
rect 65452 35848 65492 35888
rect 66796 35848 66836 35888
rect 66988 35848 67028 35888
rect 67084 35848 67124 35888
rect 67276 35848 67316 35888
rect 67372 35848 67412 35888
rect 67468 35848 67508 35888
rect 69676 35848 69716 35888
rect 69868 35848 69908 35888
rect 69964 35848 70004 35888
rect 71884 35848 71924 35888
rect 72076 35834 72116 35874
rect 72172 35848 72212 35888
rect 72748 35848 72788 35888
rect 73036 35848 73076 35888
rect 73612 35848 73652 35888
rect 73804 35848 73844 35888
rect 73996 35848 74036 35888
rect 74188 35848 74228 35888
rect 76108 35848 76148 35888
rect 76204 35848 76244 35888
rect 76300 35848 76340 35888
rect 76492 35848 76532 35888
rect 76684 35848 76724 35888
rect 76780 35848 76820 35888
rect 77068 35848 77108 35888
rect 77260 35848 77300 35888
rect 77452 35848 77492 35888
rect 77644 35848 77684 35888
rect 51340 35764 51380 35804
rect 52012 35764 52052 35804
rect 56332 35764 56372 35804
rect 61420 35764 61460 35804
rect 64204 35764 64244 35804
rect 66892 35764 66932 35804
rect 69772 35764 69812 35804
rect 73132 35764 73172 35804
rect 77164 35764 77204 35804
rect 50764 35680 50804 35720
rect 54412 35680 54452 35720
rect 56620 35680 56660 35720
rect 61804 35680 61844 35720
rect 66604 35680 66644 35720
rect 71980 35680 72020 35720
rect 76012 35680 76052 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 55180 35344 55220 35384
rect 65836 35344 65876 35384
rect 54796 35260 54836 35300
rect 55564 35260 55604 35300
rect 62668 35260 62708 35300
rect 71404 35260 71444 35300
rect 46540 35176 46580 35216
rect 46732 35176 46772 35216
rect 46828 35176 46868 35216
rect 49612 35176 49652 35216
rect 50476 35176 50516 35216
rect 50860 35176 50900 35216
rect 51340 35176 51380 35216
rect 51436 35176 51476 35216
rect 51724 35176 51764 35216
rect 52012 35176 52052 35216
rect 52108 35162 52148 35202
rect 52300 35176 52340 35216
rect 54700 35176 54740 35216
rect 54892 35176 54932 35216
rect 55084 35176 55124 35216
rect 55276 35176 55316 35216
rect 55390 35165 55430 35205
rect 55948 35176 55988 35216
rect 56812 35176 56852 35216
rect 58156 35176 58196 35216
rect 58348 35176 58388 35216
rect 58444 35176 58484 35216
rect 59788 35176 59828 35216
rect 60172 35176 60212 35216
rect 61036 35176 61076 35216
rect 62764 35176 62804 35216
rect 63052 35176 63092 35216
rect 65932 35176 65972 35216
rect 66028 35176 66068 35216
rect 66124 35176 66164 35216
rect 66412 35176 66452 35216
rect 66700 35176 66740 35216
rect 66796 35176 66836 35216
rect 67468 35176 67508 35216
rect 67852 35176 67892 35216
rect 68716 35176 68756 35216
rect 70444 35176 70484 35216
rect 70540 35176 70580 35216
rect 70636 35176 70676 35216
rect 70732 35176 70772 35216
rect 71020 35176 71060 35216
rect 71308 35176 71348 35216
rect 71884 35176 71924 35216
rect 72076 35176 72116 35216
rect 72172 35176 72212 35216
rect 72364 35176 72404 35216
rect 72556 35176 72596 35216
rect 74188 35176 74228 35216
rect 74572 35176 74612 35216
rect 75436 35176 75476 35216
rect 77068 35176 77108 35216
rect 77452 35176 77492 35216
rect 78316 35176 78356 35216
rect 51052 35008 51092 35048
rect 52492 35008 52532 35048
rect 58636 35008 58676 35048
rect 63532 35008 63572 35048
rect 64684 35008 64724 35048
rect 67084 35008 67124 35048
rect 71692 35008 71732 35048
rect 72748 35008 72788 35048
rect 46540 34924 46580 34964
rect 48460 34924 48500 34964
rect 52300 34924 52340 34964
rect 57964 34924 58004 34964
rect 58156 34924 58196 34964
rect 62188 34924 62228 34964
rect 62380 34924 62420 34964
rect 69868 34924 69908 34964
rect 71884 34924 71924 34964
rect 72460 34924 72500 34964
rect 76588 34924 76628 34964
rect 79468 34924 79508 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 50956 34588 50996 34628
rect 55564 34588 55604 34628
rect 66988 34588 67028 34628
rect 68908 34588 68948 34628
rect 77260 34588 77300 34628
rect 45964 34504 46004 34544
rect 49228 34504 49268 34544
rect 51724 34504 51764 34544
rect 52204 34504 52244 34544
rect 52684 34504 52724 34544
rect 56524 34504 56564 34544
rect 57772 34504 57812 34544
rect 61900 34504 61940 34544
rect 66604 34504 66644 34544
rect 67948 34504 67988 34544
rect 71980 34504 72020 34544
rect 77452 34504 77492 34544
rect 78028 34504 78068 34544
rect 46156 34336 46196 34376
rect 46540 34336 46580 34376
rect 47404 34336 47444 34376
rect 49228 34336 49268 34376
rect 49420 34336 49460 34376
rect 49516 34336 49556 34376
rect 50476 34336 50516 34376
rect 50572 34336 50612 34376
rect 50668 34336 50708 34376
rect 50764 34336 50804 34376
rect 50956 34336 50996 34376
rect 51148 34336 51188 34376
rect 51244 34336 51284 34376
rect 51628 34336 51668 34376
rect 51820 34336 51860 34376
rect 52204 34336 52244 34376
rect 52396 34336 52436 34376
rect 52492 34336 52532 34376
rect 53932 34336 53972 34376
rect 54124 34336 54164 34376
rect 54220 34336 54260 34376
rect 54988 34336 55028 34376
rect 55180 34336 55220 34376
rect 55852 34336 55892 34376
rect 55948 34336 55988 34376
rect 56236 34336 56276 34376
rect 57484 34336 57524 34376
rect 57580 34336 57620 34376
rect 57772 34336 57812 34376
rect 57964 34336 58004 34376
rect 58348 34336 58388 34376
rect 59212 34336 59252 34376
rect 61900 34336 61940 34376
rect 62092 34336 62132 34376
rect 62188 34336 62228 34376
rect 62572 34336 62612 34376
rect 62764 34336 62804 34376
rect 62860 34336 62900 34376
rect 63436 34336 63476 34376
rect 64300 34336 64340 34376
rect 66124 34336 66164 34376
rect 66316 34336 66356 34376
rect 66412 34336 66452 34376
rect 66988 34336 67028 34376
rect 67180 34336 67220 34376
rect 67276 34336 67316 34376
rect 67468 34336 67508 34376
rect 67564 34336 67604 34376
rect 67669 34336 67709 34376
rect 70060 34336 70100 34376
rect 70924 34336 70964 34376
rect 71308 34336 71348 34376
rect 71692 34336 71732 34376
rect 71788 34336 71828 34376
rect 71980 34336 72020 34376
rect 72172 34336 72212 34376
rect 72556 34336 72596 34376
rect 73453 34336 73493 34376
rect 76012 34336 76052 34376
rect 76204 34336 76244 34376
rect 76300 34336 76340 34376
rect 76588 34336 76628 34376
rect 76876 34336 76916 34376
rect 76972 34336 77012 34376
rect 77452 34336 77492 34376
rect 77644 34336 77684 34376
rect 77740 34336 77780 34376
rect 77932 34336 77972 34376
rect 78124 34336 78164 34376
rect 55084 34252 55124 34292
rect 62668 34252 62708 34292
rect 63052 34252 63092 34292
rect 76108 34252 76148 34292
rect 48556 34168 48596 34208
rect 54028 34168 54068 34208
rect 60364 34168 60404 34208
rect 65452 34168 65492 34208
rect 66220 34168 66260 34208
rect 74572 34168 74612 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 46444 33832 46484 33872
rect 58348 33832 58388 33872
rect 76780 33832 76820 33872
rect 52204 33748 52244 33788
rect 55276 33748 55316 33788
rect 62284 33748 62324 33788
rect 62764 33748 62804 33788
rect 63148 33748 63188 33788
rect 71692 33748 71732 33788
rect 46540 33664 46580 33704
rect 46636 33664 46676 33704
rect 46732 33664 46772 33704
rect 48940 33664 48980 33704
rect 49132 33664 49172 33704
rect 49228 33664 49268 33704
rect 52588 33664 52628 33704
rect 53452 33664 53492 33704
rect 54892 33664 54932 33704
rect 55180 33664 55220 33704
rect 58444 33664 58484 33704
rect 58540 33664 58580 33704
rect 58828 33664 58868 33704
rect 59020 33664 59060 33704
rect 54604 33580 54644 33620
rect 58636 33619 58676 33659
rect 62188 33664 62228 33704
rect 62380 33664 62420 33704
rect 62476 33664 62516 33704
rect 62668 33664 62708 33704
rect 62860 33664 62900 33704
rect 63052 33664 63092 33704
rect 63244 33664 63284 33704
rect 66220 33664 66260 33704
rect 66604 33664 66644 33704
rect 67468 33664 67508 33704
rect 71596 33664 71636 33704
rect 71788 33664 71828 33704
rect 71980 33664 72020 33704
rect 72172 33664 72212 33704
rect 72268 33664 72308 33704
rect 72460 33664 72500 33704
rect 72652 33664 72692 33704
rect 75724 33664 75764 33704
rect 75820 33664 75860 33704
rect 76012 33664 76052 33704
rect 76204 33664 76244 33704
rect 76300 33664 76340 33704
rect 76396 33664 76436 33704
rect 76492 33664 76532 33704
rect 76684 33664 76724 33704
rect 76876 33664 76916 33704
rect 76972 33664 77012 33704
rect 77260 33664 77300 33704
rect 77452 33664 77492 33704
rect 77548 33664 77588 33704
rect 72556 33580 72596 33620
rect 46252 33496 46292 33536
rect 55564 33496 55604 33536
rect 56140 33496 56180 33536
rect 59212 33496 59252 33536
rect 63724 33496 63764 33536
rect 69772 33496 69812 33536
rect 75052 33496 75092 33536
rect 77836 33496 77876 33536
rect 48940 33412 48980 33452
rect 58924 33412 58964 33452
rect 68620 33412 68660 33452
rect 71980 33412 72020 33452
rect 76012 33412 76052 33452
rect 77260 33412 77300 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 42988 33076 43028 33116
rect 47596 33076 47636 33116
rect 66508 33076 66548 33116
rect 77164 33076 77204 33116
rect 43948 32992 43988 33032
rect 46924 32992 46964 33032
rect 48076 32992 48116 33032
rect 51628 32992 51668 33032
rect 55468 32992 55508 33032
rect 61324 32992 61364 33032
rect 78124 32992 78164 33032
rect 78412 32992 78452 33032
rect 42796 32908 42836 32948
rect 45676 32824 45716 32864
rect 45868 32824 45908 32864
rect 45964 32824 46004 32864
rect 46252 32824 46292 32864
rect 46540 32824 46580 32864
rect 46636 32824 46676 32864
rect 47116 32824 47156 32864
rect 47308 32824 47348 32864
rect 47500 32824 47540 32864
rect 47692 32824 47732 32864
rect 48268 32824 48308 32864
rect 48652 32824 48692 32864
rect 49516 32824 49556 32864
rect 50860 32824 50900 32864
rect 51052 32824 51092 32864
rect 51244 32824 51284 32864
rect 51436 32824 51476 32864
rect 53644 32824 53684 32864
rect 53740 32824 53780 32864
rect 53836 32824 53876 32864
rect 53932 32824 53972 32864
rect 54796 32824 54836 32864
rect 54892 32824 54932 32864
rect 54988 32824 55028 32864
rect 55180 32824 55220 32864
rect 55276 32824 55316 32864
rect 55468 32824 55508 32864
rect 55660 32824 55700 32864
rect 56044 32824 56084 32864
rect 56908 32824 56948 32864
rect 58252 32824 58292 32864
rect 58444 32824 58484 32864
rect 58540 32824 58580 32864
rect 59116 32824 59156 32864
rect 59980 32824 60020 32864
rect 62476 32824 62516 32864
rect 62572 32824 62612 32864
rect 62668 32824 62708 32864
rect 63628 32824 63668 32864
rect 64492 32824 64532 32864
rect 66028 32824 66068 32864
rect 66124 32824 66164 32864
rect 66220 32824 66260 32864
rect 66316 32824 66356 32864
rect 66508 32824 66548 32864
rect 66700 32824 66740 32864
rect 66796 32824 66836 32864
rect 68812 32824 68852 32864
rect 68908 32824 68948 32864
rect 69100 32824 69140 32864
rect 69676 32824 69716 32864
rect 70540 32824 70580 32864
rect 72172 32824 72212 32864
rect 72556 32824 72596 32864
rect 73420 32813 73460 32853
rect 74764 32824 74804 32864
rect 75148 32824 75188 32864
rect 76012 32824 76052 32864
rect 77452 32824 77492 32864
rect 77740 32824 77780 32864
rect 77836 32824 77876 32864
rect 78316 32824 78356 32864
rect 78508 32824 78548 32864
rect 47212 32740 47252 32780
rect 50956 32740 50996 32780
rect 51340 32740 51380 32780
rect 58348 32740 58388 32780
rect 58732 32740 58772 32780
rect 63244 32740 63284 32780
rect 69292 32740 69332 32780
rect 45772 32656 45812 32696
rect 50668 32656 50708 32696
rect 58060 32656 58100 32696
rect 61132 32656 61172 32696
rect 62380 32656 62420 32696
rect 65644 32656 65684 32696
rect 69004 32656 69044 32696
rect 71692 32656 71732 32696
rect 74572 32656 74612 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 48268 32320 48308 32360
rect 48748 32320 48788 32360
rect 54220 32320 54260 32360
rect 62764 32320 62804 32360
rect 69964 32320 70004 32360
rect 75916 32320 75956 32360
rect 45868 32236 45908 32276
rect 58732 32236 58772 32276
rect 63436 32236 63476 32276
rect 66028 32236 66068 32276
rect 71980 32236 72020 32276
rect 76780 32236 76820 32276
rect 77068 32236 77108 32276
rect 42412 32152 42452 32192
rect 42508 32152 42548 32192
rect 42604 32152 42644 32192
rect 42700 32152 42740 32192
rect 42892 32152 42932 32192
rect 43084 32152 43124 32192
rect 43276 32152 43316 32192
rect 43660 32152 43700 32192
rect 44524 32152 44564 32192
rect 46252 32152 46292 32192
rect 47116 32152 47156 32192
rect 48460 32152 48500 32192
rect 48844 32152 48884 32192
rect 48940 32152 48980 32192
rect 49036 32107 49076 32147
rect 49420 32152 49460 32192
rect 51148 32152 51188 32192
rect 51532 32152 51572 32192
rect 52396 32152 52436 32192
rect 54124 32152 54164 32192
rect 54316 32152 54356 32192
rect 54412 32152 54452 32192
rect 54604 32152 54644 32192
rect 54700 32152 54740 32192
rect 54796 32152 54836 32192
rect 54892 32152 54932 32192
rect 58348 32152 58388 32192
rect 58636 32152 58676 32192
rect 59212 32152 59252 32192
rect 59404 32152 59444 32192
rect 59596 32152 59636 32192
rect 59692 32152 59732 32192
rect 59884 32152 59924 32192
rect 60364 32152 60404 32192
rect 60748 32152 60788 32192
rect 61612 32152 61652 32192
rect 63052 32152 63092 32192
rect 63340 32179 63380 32219
rect 63916 32152 63956 32192
rect 64108 32173 64148 32213
rect 64300 32152 64340 32192
rect 64492 32152 64532 32192
rect 65356 32152 65396 32192
rect 65548 32152 65588 32192
rect 66124 32152 66164 32192
rect 66412 32152 66452 32192
rect 66700 32152 66740 32192
rect 67084 32152 67124 32192
rect 67948 32152 67988 32192
rect 69772 32152 69812 32192
rect 69868 32152 69908 32192
rect 70060 32152 70100 32192
rect 70252 32152 70292 32192
rect 70348 32152 70388 32192
rect 70444 32152 70484 32192
rect 70540 32152 70580 32192
rect 70828 32152 70868 32192
rect 70924 32152 70964 32192
rect 71116 32152 71156 32192
rect 71596 32152 71636 32192
rect 71884 32152 71924 32192
rect 72460 32152 72500 32192
rect 72652 32152 72692 32192
rect 75820 32152 75860 32192
rect 76012 32152 76052 32192
rect 76108 32152 76148 32192
rect 76684 32152 76724 32192
rect 76876 32152 76916 32192
rect 77452 32152 77492 32192
rect 78316 32152 78356 32192
rect 59308 32068 59348 32108
rect 79468 32068 79508 32108
rect 40588 31984 40628 32024
rect 53548 31984 53588 32024
rect 56620 31984 56660 32024
rect 59020 31984 59060 32024
rect 63724 31984 63764 32024
rect 65452 31984 65492 32024
rect 65740 31984 65780 32024
rect 72268 31984 72308 32024
rect 72556 31984 72596 32024
rect 72844 31984 72884 32024
rect 74092 31984 74132 32024
rect 42988 31900 43028 31940
rect 45676 31900 45716 31940
rect 49612 31900 49652 31940
rect 59884 31900 59924 31940
rect 64012 31900 64052 31940
rect 64396 31900 64436 31940
rect 69100 31900 69140 31940
rect 71116 31900 71156 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 42700 31564 42740 31604
rect 43948 31564 43988 31604
rect 48844 31564 48884 31604
rect 51148 31564 51188 31604
rect 51820 31564 51860 31604
rect 55180 31564 55220 31604
rect 63052 31564 63092 31604
rect 66412 31564 66452 31604
rect 71116 31564 71156 31604
rect 76012 31564 76052 31604
rect 48364 31480 48404 31520
rect 49708 31480 49748 31520
rect 61132 31480 61172 31520
rect 50956 31438 50996 31478
rect 63628 31480 63668 31520
rect 67276 31480 67316 31520
rect 68812 31480 68852 31520
rect 72268 31480 72308 31520
rect 77836 31480 77876 31520
rect 51628 31396 51668 31436
rect 60652 31396 60692 31436
rect 70924 31396 70964 31436
rect 40492 31312 40532 31352
rect 41356 31312 41396 31352
rect 43084 31312 43124 31352
rect 43372 31312 43412 31352
rect 43660 31312 43700 31352
rect 43756 31312 43796 31352
rect 43948 31312 43988 31352
rect 48556 31312 48596 31352
rect 48652 31312 48692 31352
rect 48844 31312 48884 31352
rect 49228 31312 49268 31352
rect 49420 31312 49460 31352
rect 49516 31312 49556 31352
rect 49708 31312 49748 31352
rect 49900 31312 49940 31352
rect 49996 31312 50036 31352
rect 50284 31312 50324 31352
rect 50572 31312 50612 31352
rect 50668 31312 50708 31352
rect 51148 31312 51188 31352
rect 51340 31312 51380 31352
rect 51436 31312 51476 31352
rect 53164 31312 53204 31352
rect 54028 31312 54068 31352
rect 55564 31312 55604 31352
rect 55756 31312 55796 31352
rect 56524 31312 56564 31352
rect 57388 31312 57428 31352
rect 59596 31312 59636 31352
rect 59788 31312 59828 31352
rect 59884 31312 59924 31352
rect 62572 31312 62612 31352
rect 62764 31312 62804 31352
rect 62860 31312 62900 31352
rect 63052 31312 63092 31352
rect 63244 31312 63284 31352
rect 63358 31323 63398 31363
rect 66412 31312 66452 31352
rect 66604 31312 66644 31352
rect 66700 31312 66740 31352
rect 66892 31312 66932 31352
rect 67084 31312 67124 31352
rect 70540 31312 70580 31352
rect 70636 31312 70676 31352
rect 70732 31312 70772 31352
rect 71404 31312 71444 31352
rect 71596 31312 71636 31352
rect 73996 31312 74036 31352
rect 74860 31312 74900 31352
rect 76972 31312 77012 31352
rect 77164 31312 77204 31352
rect 77452 31312 77492 31352
rect 77644 31312 77684 31352
rect 40108 31228 40148 31268
rect 42988 31228 43028 31268
rect 52780 31228 52820 31268
rect 55660 31228 55700 31268
rect 56140 31228 56180 31268
rect 62668 31228 62708 31268
rect 66988 31228 67028 31268
rect 71500 31228 71540 31268
rect 73612 31228 73652 31268
rect 77068 31228 77108 31268
rect 77548 31228 77588 31268
rect 42508 31144 42548 31184
rect 49324 31144 49364 31184
rect 51820 31144 51860 31184
rect 55180 31144 55220 31184
rect 58540 31144 58580 31184
rect 59692 31144 59732 31184
rect 60460 31144 60500 31184
rect 70444 31144 70484 31184
rect 71116 31144 71156 31184
rect 76012 31144 76052 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 40972 30808 41012 30848
rect 52108 30808 52148 30848
rect 56044 30808 56084 30848
rect 60940 30808 60980 30848
rect 61708 30808 61748 30848
rect 62764 30808 62804 30848
rect 75436 30808 75476 30848
rect 43372 30724 43412 30764
rect 48076 30724 48116 30764
rect 50860 30724 50900 30764
rect 55468 30724 55508 30764
rect 57772 30724 57812 30764
rect 71308 30724 71348 30764
rect 74860 30724 74900 30764
rect 42796 30629 42836 30669
rect 42988 30640 43028 30680
rect 43084 30640 43124 30680
rect 43276 30640 43316 30680
rect 43468 30640 43508 30680
rect 43948 30640 43988 30680
rect 44140 30640 44180 30680
rect 44236 30640 44276 30680
rect 44908 30640 44948 30680
rect 45004 30640 45044 30680
rect 45100 30640 45140 30680
rect 45196 30640 45236 30680
rect 45868 30640 45908 30680
rect 46060 30640 46100 30680
rect 46252 30640 46292 30680
rect 46348 30640 46388 30680
rect 46540 30640 46580 30680
rect 48460 30640 48500 30680
rect 49324 30640 49364 30680
rect 50764 30640 50804 30680
rect 50956 30640 50996 30680
rect 51148 30640 51188 30680
rect 51340 30640 51380 30680
rect 54508 30640 54548 30680
rect 54700 30640 54740 30680
rect 54796 30640 54836 30680
rect 55084 30640 55124 30680
rect 55372 30640 55412 30680
rect 55948 30640 55988 30680
rect 56140 30640 56180 30680
rect 56236 30640 56276 30680
rect 56428 30640 56468 30680
rect 56620 30640 56660 30680
rect 58156 30640 58196 30680
rect 59020 30651 59060 30691
rect 61132 30640 61172 30680
rect 61324 30640 61364 30680
rect 62668 30640 62708 30680
rect 62860 30640 62900 30680
rect 62956 30640 62996 30680
rect 63148 30640 63188 30680
rect 63532 30640 63572 30680
rect 64396 30640 64436 30680
rect 65932 30640 65972 30680
rect 66124 30653 66164 30693
rect 68236 30640 68276 30680
rect 68620 30640 68660 30680
rect 69484 30640 69524 30680
rect 70924 30640 70964 30680
rect 71212 30640 71252 30680
rect 71788 30640 71828 30680
rect 72172 30640 72212 30680
rect 73036 30640 73076 30680
rect 74956 30640 74996 30680
rect 75052 30640 75092 30680
rect 75148 30640 75188 30680
rect 75340 30640 75380 30680
rect 75532 30640 75572 30680
rect 75628 30640 75668 30680
rect 76204 30640 76244 30680
rect 76492 30640 76532 30680
rect 76588 30640 76628 30680
rect 77068 30640 77108 30680
rect 77452 30640 77492 30680
rect 78316 30640 78356 30680
rect 40588 30556 40628 30596
rect 41164 30556 41204 30596
rect 42412 30556 42452 30596
rect 51532 30556 51572 30596
rect 51916 30556 51956 30596
rect 43948 30472 43988 30512
rect 44428 30472 44468 30512
rect 47020 30472 47060 30512
rect 52300 30472 52340 30512
rect 53260 30514 53300 30554
rect 56524 30556 56564 30596
rect 60556 30556 60596 30596
rect 60748 30556 60788 30596
rect 61516 30556 61556 30596
rect 54508 30472 54548 30512
rect 55756 30472 55796 30512
rect 66508 30472 66548 30512
rect 71596 30472 71636 30512
rect 76876 30472 76916 30512
rect 79468 30472 79508 30512
rect 40780 30388 40820 30428
rect 40972 30388 41012 30428
rect 42604 30388 42644 30428
rect 42796 30388 42836 30428
rect 45964 30388 46004 30428
rect 46540 30388 46580 30428
rect 50476 30388 50516 30428
rect 51244 30388 51284 30428
rect 51724 30388 51764 30428
rect 52108 30388 52148 30428
rect 60172 30388 60212 30428
rect 60364 30388 60404 30428
rect 60940 30388 60980 30428
rect 61228 30388 61268 30428
rect 61708 30388 61748 30428
rect 65548 30388 65588 30428
rect 66028 30388 66068 30428
rect 70636 30388 70676 30428
rect 74188 30388 74228 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 40588 30052 40628 30092
rect 45964 30052 46004 30092
rect 46252 30052 46292 30092
rect 50956 30052 50996 30092
rect 54796 30052 54836 30092
rect 56428 30052 56468 30092
rect 58828 30052 58868 30092
rect 63724 30052 63764 30092
rect 69100 30052 69140 30092
rect 69676 30052 69716 30092
rect 71500 30052 71540 30092
rect 75724 30052 75764 30092
rect 77068 30052 77108 30092
rect 38956 29968 38996 30008
rect 42316 29968 42356 30008
rect 55756 29968 55796 30008
rect 56620 29968 56660 30008
rect 58252 29968 58292 30008
rect 60460 29968 60500 30008
rect 65068 29968 65108 30008
rect 70348 29968 70388 30008
rect 73900 29968 73940 30008
rect 76588 29968 76628 30008
rect 77548 29968 77588 30008
rect 40012 29884 40052 29924
rect 40396 29884 40436 29924
rect 42124 29884 42164 29924
rect 49324 29884 49364 29924
rect 56236 29884 56276 29924
rect 59020 29871 59060 29911
rect 69292 29884 69332 29924
rect 69484 29884 69524 29924
rect 75052 29884 75092 29924
rect 40780 29800 40820 29840
rect 40876 29800 40916 29840
rect 40972 29800 41012 29840
rect 41260 29800 41300 29840
rect 41452 29800 41492 29840
rect 41644 29800 41684 29840
rect 41836 29800 41876 29840
rect 41932 29800 41972 29840
rect 43948 29800 43988 29840
rect 44812 29800 44852 29840
rect 46156 29800 46196 29840
rect 46348 29800 46388 29840
rect 46540 29800 46580 29840
rect 46924 29800 46964 29840
rect 47788 29800 47828 29840
rect 49708 29800 49748 29840
rect 49804 29800 49844 29840
rect 49900 29779 49940 29819
rect 49996 29800 50036 29840
rect 50284 29800 50324 29840
rect 50572 29800 50612 29840
rect 50668 29800 50708 29840
rect 51628 29800 51668 29840
rect 52492 29800 52532 29840
rect 54796 29800 54836 29840
rect 54988 29800 55028 29840
rect 55084 29800 55124 29840
rect 55660 29800 55700 29840
rect 55852 29800 55892 29840
rect 59212 29800 59252 29840
rect 59308 29800 59348 29840
rect 59404 29800 59444 29840
rect 59500 29800 59540 29840
rect 59788 29800 59828 29840
rect 60076 29800 60116 29840
rect 60172 29800 60212 29840
rect 61036 29800 61076 29840
rect 61900 29800 61940 29840
rect 63340 29842 63380 29882
rect 63244 29800 63284 29840
rect 63436 29800 63476 29840
rect 63532 29800 63572 29840
rect 63724 29800 63764 29840
rect 63916 29800 63956 29840
rect 64012 29800 64052 29840
rect 64684 29800 64724 29840
rect 64876 29800 64916 29840
rect 65356 29800 65396 29840
rect 65452 29800 65492 29840
rect 65740 29800 65780 29840
rect 66412 29800 66452 29840
rect 67276 29800 67316 29840
rect 69868 29800 69908 29840
rect 70060 29800 70100 29840
rect 70156 29800 70196 29840
rect 70348 29800 70388 29840
rect 70540 29800 70580 29840
rect 70636 29800 70676 29840
rect 70828 29800 70868 29840
rect 71020 29800 71060 29840
rect 71116 29800 71156 29840
rect 71500 29800 71540 29840
rect 71692 29800 71732 29840
rect 71788 29800 71828 29840
rect 71980 29800 72020 29840
rect 72076 29800 72116 29840
rect 72172 29800 72212 29840
rect 75340 29800 75380 29840
rect 75436 29800 75476 29840
rect 75532 29800 75572 29840
rect 75724 29800 75764 29840
rect 76012 29800 76052 29840
rect 76492 29800 76532 29840
rect 76684 29800 76724 29840
rect 41356 29716 41396 29756
rect 43564 29716 43604 29756
rect 51244 29716 51284 29756
rect 60652 29716 60692 29756
rect 64780 29716 64820 29756
rect 66028 29716 66068 29756
rect 70924 29716 70964 29756
rect 75916 29758 75956 29798
rect 77068 29800 77108 29840
rect 77260 29800 77300 29840
rect 77356 29800 77396 29840
rect 40204 29632 40244 29672
rect 41068 29632 41108 29672
rect 41740 29632 41780 29672
rect 45964 29632 46004 29672
rect 48940 29632 48980 29672
rect 49516 29632 49556 29672
rect 53644 29632 53684 29672
rect 63052 29632 63092 29672
rect 68428 29632 68468 29672
rect 69676 29632 69716 29672
rect 69964 29632 70004 29672
rect 74860 29632 74900 29672
rect 75244 29632 75284 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 49612 29296 49652 29336
rect 51052 29296 51092 29336
rect 55276 29296 55316 29336
rect 60460 29296 60500 29336
rect 63436 29296 63476 29336
rect 70252 29296 70292 29336
rect 70732 29296 70772 29336
rect 71692 29296 71732 29336
rect 75820 29296 75860 29336
rect 45964 29212 46004 29252
rect 60940 29212 60980 29252
rect 65740 29212 65780 29252
rect 67660 29212 67700 29252
rect 76492 29212 76532 29252
rect 38476 29128 38516 29168
rect 38860 29128 38900 29168
rect 39724 29128 39764 29168
rect 41356 29128 41396 29168
rect 41452 29128 41492 29168
rect 41740 29128 41780 29168
rect 42028 29128 42068 29168
rect 42124 29128 42164 29168
rect 42316 29128 42356 29168
rect 45100 29128 45140 29168
rect 45292 29128 45332 29168
rect 45388 29128 45428 29168
rect 46060 29128 46100 29168
rect 46348 29128 46388 29168
rect 50188 29128 50228 29168
rect 50380 29128 50420 29168
rect 50476 29128 50516 29168
rect 50860 29128 50900 29168
rect 50956 29128 50996 29168
rect 51148 29128 51188 29168
rect 52876 29128 52916 29168
rect 53260 29092 53300 29132
rect 54124 29128 54164 29168
rect 55468 29128 55508 29168
rect 55564 29128 55604 29168
rect 55660 29128 55700 29168
rect 55756 29128 55796 29168
rect 56140 29128 56180 29168
rect 56524 29128 56564 29168
rect 57388 29128 57428 29168
rect 59596 29128 59636 29168
rect 59692 29128 59732 29168
rect 59884 29128 59924 29168
rect 60364 29128 60404 29168
rect 60556 29128 60596 29168
rect 60652 29128 60692 29168
rect 60844 29128 60884 29168
rect 61036 29128 61076 29168
rect 63340 29117 63380 29157
rect 63532 29128 63572 29168
rect 63628 29128 63668 29168
rect 63820 29128 63860 29168
rect 63916 29128 63956 29168
rect 64012 29128 64052 29168
rect 64108 29128 64148 29168
rect 65644 29128 65684 29168
rect 65836 29128 65876 29168
rect 65932 29128 65972 29168
rect 68044 29128 68084 29168
rect 68908 29128 68948 29168
rect 70348 29128 70388 29168
rect 70444 29128 70484 29168
rect 70540 29128 70580 29168
rect 73804 29128 73844 29168
rect 74668 29128 74708 29168
rect 76108 29128 76148 29168
rect 76396 29128 76436 29168
rect 49420 29044 49460 29084
rect 49996 29044 50036 29084
rect 59212 29044 59252 29084
rect 73420 29086 73460 29126
rect 77068 29128 77108 29168
rect 77452 29128 77492 29168
rect 78316 29128 78356 29168
rect 70060 29044 70100 29084
rect 70924 29044 70964 29084
rect 71116 29044 71156 29084
rect 71500 29044 71540 29084
rect 72076 29044 72116 29084
rect 41068 28960 41108 29000
rect 42508 28960 42548 29000
rect 44716 28960 44756 29000
rect 45100 28960 45140 29000
rect 45676 28960 45716 29000
rect 49804 28960 49844 29000
rect 59404 28960 59444 29000
rect 62380 28960 62420 29000
rect 67468 28960 67508 29000
rect 71308 28960 71348 29000
rect 76780 28960 76820 29000
rect 40876 28876 40916 28916
rect 42316 28876 42356 28916
rect 50188 28876 50228 28916
rect 58540 28876 58580 28916
rect 59884 28876 59924 28916
rect 71884 28876 71924 28916
rect 79468 28876 79508 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 41068 28540 41108 28580
rect 41644 28540 41684 28580
rect 44620 28540 44660 28580
rect 51340 28540 51380 28580
rect 54604 28540 54644 28580
rect 56044 28540 56084 28580
rect 56236 28540 56276 28580
rect 61036 28540 61076 28580
rect 61612 28540 61652 28580
rect 76780 28540 76820 28580
rect 47596 28456 47636 28496
rect 49324 28456 49364 28496
rect 51724 28456 51764 28496
rect 52300 28456 52340 28496
rect 52492 28456 52532 28496
rect 57772 28456 57812 28496
rect 64492 28456 64532 28496
rect 70924 28456 70964 28496
rect 39532 28372 39572 28412
rect 40108 28372 40148 28412
rect 46252 28372 46292 28412
rect 51148 28372 51188 28412
rect 58924 28372 58964 28412
rect 59596 28372 59636 28412
rect 61228 28372 61268 28412
rect 61420 28372 61460 28412
rect 73804 28372 73844 28412
rect 40300 28288 40340 28328
rect 40492 28288 40532 28328
rect 40588 28288 40628 28328
rect 41068 28288 41108 28328
rect 41260 28288 41300 28328
rect 41356 28288 41396 28328
rect 41548 28288 41588 28328
rect 41740 28288 41780 28328
rect 41932 28288 41972 28328
rect 42316 28288 42356 28328
rect 43213 28288 43253 28328
rect 44620 28288 44660 28328
rect 44812 28288 44852 28328
rect 44908 28288 44948 28328
rect 45100 28288 45140 28328
rect 45196 28288 45236 28328
rect 45292 28288 45332 28328
rect 45388 28288 45428 28328
rect 45580 28288 45620 28328
rect 45772 28288 45812 28328
rect 45868 28288 45908 28328
rect 46636 28288 46676 28328
rect 46828 28288 46868 28328
rect 49996 28288 50036 28328
rect 50188 28288 50228 28328
rect 50284 28288 50324 28328
rect 50476 28288 50516 28328
rect 50572 28288 50612 28328
rect 50668 28288 50708 28328
rect 50764 28288 50804 28328
rect 51628 28288 51668 28328
rect 51820 28288 51860 28328
rect 52972 28288 53012 28328
rect 55372 28288 55412 28328
rect 55660 28288 55700 28328
rect 55756 28288 55796 28328
rect 56236 28288 56276 28328
rect 56428 28288 56468 28328
rect 56524 28288 56564 28328
rect 56716 28288 56756 28328
rect 56908 28288 56948 28328
rect 59116 28288 59156 28328
rect 59212 28288 59252 28328
rect 59308 28288 59348 28328
rect 60172 28288 60212 28328
rect 60364 28288 60404 28328
rect 60460 28288 60500 28328
rect 60652 28288 60692 28328
rect 60748 28288 60788 28328
rect 60844 28288 60884 28328
rect 62284 28288 62324 28328
rect 63148 28288 63188 28328
rect 64780 28288 64820 28328
rect 64876 28288 64916 28328
rect 65164 28288 65204 28328
rect 66124 28288 66164 28328
rect 66988 28288 67028 28328
rect 70252 28288 70292 28328
rect 70540 28288 70580 28328
rect 70636 28288 70676 28328
rect 71788 28288 71828 28328
rect 72652 28288 72692 28328
rect 75244 28288 75284 28328
rect 75436 28288 75476 28328
rect 75532 28288 75572 28328
rect 76780 28288 76820 28328
rect 76972 28288 77012 28328
rect 77068 28288 77108 28328
rect 77260 28288 77300 28328
rect 77452 28288 77492 28328
rect 46732 28204 46772 28244
rect 56812 28204 56852 28244
rect 61900 28204 61940 28244
rect 65740 28204 65780 28244
rect 71404 28204 71444 28244
rect 75340 28204 75380 28244
rect 77356 28204 77396 28244
rect 39724 28120 39764 28160
rect 39916 28120 39956 28160
rect 40396 28120 40436 28160
rect 44332 28120 44372 28160
rect 45676 28120 45716 28160
rect 46060 28120 46100 28160
rect 50092 28120 50132 28160
rect 58732 28120 58772 28160
rect 59404 28120 59444 28160
rect 59788 28120 59828 28160
rect 60268 28120 60308 28160
rect 61036 28120 61076 28160
rect 64300 28120 64340 28160
rect 68140 28120 68180 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 3820 27784 3860 27824
rect 41452 27784 41492 27824
rect 43564 27784 43604 27824
rect 51244 27784 51284 27824
rect 59692 27784 59732 27824
rect 63916 27784 63956 27824
rect 71116 27784 71156 27824
rect 37804 27700 37844 27740
rect 40492 27700 40532 27740
rect 45964 27700 46004 27740
rect 46636 27700 46676 27740
rect 47692 27700 47732 27740
rect 48844 27700 48884 27740
rect 51628 27700 51668 27740
rect 52012 27700 52052 27740
rect 57292 27700 57332 27740
rect 59980 27700 60020 27740
rect 60556 27700 60596 27740
rect 70732 27700 70772 27740
rect 3724 27616 3764 27656
rect 38188 27616 38228 27656
rect 39052 27616 39092 27656
rect 40396 27616 40436 27656
rect 40588 27616 40628 27656
rect 40684 27616 40724 27656
rect 41068 27616 41108 27656
rect 41260 27616 41300 27656
rect 44716 27616 44756 27656
rect 45580 27616 45620 27656
rect 46252 27616 46292 27656
rect 46540 27616 46580 27656
rect 47116 27616 47156 27656
rect 47308 27616 47348 27656
rect 47404 27616 47444 27656
rect 47596 27616 47636 27656
rect 47788 27616 47828 27656
rect 47980 27616 48020 27656
rect 49228 27616 49268 27656
rect 50092 27616 50132 27656
rect 51532 27616 51572 27656
rect 51724 27616 51764 27656
rect 51820 27616 51860 27656
rect 52396 27616 52436 27656
rect 53293 27616 53333 27656
rect 54604 27616 54644 27656
rect 54796 27616 54836 27656
rect 54892 27616 54932 27656
rect 55180 27616 55220 27656
rect 55372 27616 55412 27656
rect 55468 27616 55508 27656
rect 55660 27616 55700 27656
rect 55756 27616 55796 27656
rect 55852 27616 55892 27656
rect 55948 27616 55988 27656
rect 57676 27616 57716 27656
rect 58540 27616 58580 27656
rect 59884 27616 59924 27656
rect 60076 27616 60116 27656
rect 60172 27616 60212 27656
rect 60940 27616 60980 27656
rect 61804 27616 61844 27656
rect 63724 27616 63764 27656
rect 63820 27616 63860 27656
rect 64012 27616 64052 27656
rect 64780 27616 64820 27656
rect 64876 27616 64916 27656
rect 64972 27616 65012 27656
rect 65164 27616 65204 27656
rect 65356 27616 65396 27656
rect 65452 27616 65492 27656
rect 65644 27616 65684 27656
rect 65836 27616 65876 27656
rect 69580 27616 69620 27656
rect 69772 27616 69812 27656
rect 69868 27616 69908 27656
rect 70060 27616 70100 27656
rect 70252 27616 70292 27656
rect 70348 27616 70388 27656
rect 70636 27616 70676 27656
rect 70828 27616 70868 27656
rect 71020 27616 71060 27656
rect 71212 27616 71252 27656
rect 71308 27616 71348 27656
rect 71500 27616 71540 27656
rect 71692 27629 71732 27669
rect 74860 27616 74900 27656
rect 75052 27616 75092 27656
rect 75148 27616 75188 27656
rect 75436 27616 75476 27656
rect 75628 27616 75668 27656
rect 75724 27616 75764 27656
rect 76684 27616 76724 27656
rect 76780 27616 76820 27656
rect 76876 27616 76916 27656
rect 77164 27616 77204 27656
rect 77356 27616 77396 27656
rect 41644 27532 41684 27572
rect 65740 27532 65780 27572
rect 67564 27532 67604 27572
rect 46924 27448 46964 27488
rect 54604 27448 54644 27488
rect 56140 27448 56180 27488
rect 59692 27448 59732 27488
rect 65164 27448 65204 27488
rect 66220 27448 66260 27488
rect 69388 27448 69428 27488
rect 69580 27448 69620 27488
rect 70060 27448 70100 27488
rect 71884 27448 71924 27488
rect 73516 27448 73556 27488
rect 77548 27448 77588 27488
rect 3820 27364 3860 27404
rect 40204 27364 40244 27404
rect 41164 27364 41204 27404
rect 41452 27364 41492 27404
rect 47116 27364 47156 27404
rect 51244 27364 51284 27404
rect 54412 27364 54452 27404
rect 55180 27364 55220 27404
rect 62956 27364 62996 27404
rect 67372 27364 67412 27404
rect 71596 27364 71636 27404
rect 74860 27364 74900 27404
rect 75436 27364 75476 27404
rect 77260 27364 77300 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 39724 27028 39764 27068
rect 41164 27028 41204 27068
rect 49516 27028 49556 27068
rect 51820 27028 51860 27068
rect 52108 27028 52148 27068
rect 54220 27028 54260 27068
rect 58540 27028 58580 27068
rect 60172 27028 60212 27068
rect 60844 27028 60884 27068
rect 63820 27028 63860 27068
rect 68812 27028 68852 27068
rect 71980 27028 72020 27068
rect 72172 27028 72212 27068
rect 76876 27028 76916 27068
rect 35116 26944 35156 26984
rect 38284 26944 38324 26984
rect 39340 26944 39380 26984
rect 58156 26944 58196 26984
rect 61132 26944 61172 26984
rect 62092 26944 62132 26984
rect 39148 26860 39188 26900
rect 39532 26860 39572 26900
rect 50398 26863 50438 26903
rect 57964 26860 58004 26900
rect 58348 26860 58388 26900
rect 60364 26860 60404 26900
rect 69004 26860 69044 26900
rect 71788 26860 71828 26900
rect 72364 26860 72404 26900
rect 75436 26860 75476 26900
rect 35020 26776 35060 26816
rect 35212 26776 35252 26816
rect 36076 26776 36116 26816
rect 36940 26776 36980 26816
rect 39916 26776 39956 26816
rect 40012 26776 40052 26816
rect 40108 26776 40148 26816
rect 40204 26776 40244 26816
rect 40492 26776 40532 26816
rect 40780 26776 40820 26816
rect 40876 26776 40916 26816
rect 41356 26776 41396 26816
rect 41548 26776 41588 26816
rect 42124 26776 42164 26816
rect 42988 26776 43028 26816
rect 45388 26776 45428 26816
rect 46828 26776 46868 26816
rect 47116 26776 47156 26816
rect 47500 26776 47540 26816
rect 48364 26776 48404 26816
rect 50572 26787 50612 26827
rect 50764 26776 50804 26816
rect 50860 26776 50900 26816
rect 51148 26776 51188 26816
rect 51436 26776 51476 26816
rect 51532 26776 51572 26816
rect 52012 26776 52052 26816
rect 52204 26776 52244 26816
rect 55372 26776 55412 26816
rect 56236 26776 56276 26816
rect 58828 26776 58868 26816
rect 59020 26776 59060 26816
rect 59116 26776 59156 26816
rect 59500 26776 59540 26816
rect 59788 26776 59828 26816
rect 59884 26776 59924 26816
rect 60748 26776 60788 26816
rect 60940 26776 60980 26816
rect 63820 26776 63860 26816
rect 64012 26776 64052 26816
rect 64108 26776 64148 26816
rect 66796 26776 66836 26816
rect 67660 26776 67700 26816
rect 68332 26776 68372 26816
rect 68524 26776 68564 26816
rect 68620 26776 68660 26816
rect 69196 26776 69236 26816
rect 69580 26776 69620 26816
rect 70444 26776 70484 26816
rect 73036 26776 73076 26816
rect 73420 26812 73460 26852
rect 74284 26776 74324 26816
rect 75628 26776 75668 26816
rect 75724 26776 75764 26816
rect 75820 26776 75860 26816
rect 75916 26776 75956 26816
rect 76204 26776 76244 26816
rect 76492 26776 76532 26816
rect 76588 26776 76628 26816
rect 77452 26776 77492 26816
rect 78316 26776 78356 26816
rect 35692 26692 35732 26732
rect 41452 26692 41492 26732
rect 41740 26692 41780 26732
rect 56620 26692 56660 26732
rect 68044 26692 68084 26732
rect 77068 26692 77108 26732
rect 38092 26608 38132 26648
rect 39724 26608 39764 26648
rect 44140 26608 44180 26648
rect 49516 26608 49556 26648
rect 50188 26608 50228 26648
rect 50668 26608 50708 26648
rect 58540 26608 58580 26648
rect 58924 26608 58964 26648
rect 60556 26608 60596 26648
rect 65644 26608 65684 26648
rect 68428 26608 68468 26648
rect 71596 26608 71636 26648
rect 71980 26608 72020 26648
rect 72172 26608 72212 26648
rect 79468 26608 79508 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 35692 26272 35732 26312
rect 39052 26272 39092 26312
rect 40588 26272 40628 26312
rect 40780 26272 40820 26312
rect 41548 26272 41588 26312
rect 46540 26272 46580 26312
rect 52108 26272 52148 26312
rect 56428 26272 56468 26312
rect 59020 26272 59060 26312
rect 61132 26272 61172 26312
rect 67756 26272 67796 26312
rect 69580 26272 69620 26312
rect 70636 26272 70676 26312
rect 74668 26272 74708 26312
rect 76876 26272 76916 26312
rect 35020 26188 35060 26228
rect 48844 26188 48884 26228
rect 51532 26188 51572 26228
rect 55660 26188 55700 26228
rect 61612 26188 61652 26228
rect 64780 26188 64820 26228
rect 71308 26188 71348 26228
rect 71884 26188 71924 26228
rect 75244 26188 75284 26228
rect 33148 26104 33188 26144
rect 33964 26104 34004 26144
rect 34348 26104 34388 26144
rect 34636 26104 34676 26144
rect 34924 26104 34964 26144
rect 35500 26104 35540 26144
rect 35596 26104 35636 26144
rect 35788 26104 35828 26144
rect 39244 26104 39284 26144
rect 39436 26104 39476 26144
rect 39532 26104 39572 26144
rect 39724 26104 39764 26144
rect 39916 26104 39956 26144
rect 40012 26104 40052 26144
rect 41356 26104 41396 26144
rect 41452 26104 41492 26144
rect 41644 26104 41684 26144
rect 43852 26104 43892 26144
rect 44236 26104 44276 26144
rect 45100 26104 45140 26144
rect 46444 26104 46484 26144
rect 46636 26104 46676 26144
rect 46732 26104 46772 26144
rect 47788 26104 47828 26144
rect 48652 26104 48692 26144
rect 49228 26104 49268 26144
rect 50092 26104 50132 26144
rect 51436 26104 51476 26144
rect 51628 26104 51668 26144
rect 51724 26104 51764 26144
rect 52492 26104 52532 26144
rect 52684 26104 52724 26144
rect 54988 26104 55028 26144
rect 55180 26104 55220 26144
rect 55756 26104 55796 26144
rect 56044 26104 56084 26144
rect 56332 26104 56372 26144
rect 56524 26104 56564 26144
rect 56620 26104 56660 26144
rect 56812 26104 56852 26144
rect 57004 26104 57044 26144
rect 57100 26104 57140 26144
rect 58348 26104 58388 26144
rect 58540 26104 58580 26144
rect 58636 26104 58676 26144
rect 59308 26081 59348 26121
rect 59500 26104 59540 26144
rect 59692 26104 59732 26144
rect 59788 26104 59828 26144
rect 59980 26104 60020 26144
rect 61996 26104 62036 26144
rect 62860 26104 62900 26144
rect 64204 26104 64244 26144
rect 64300 26104 64340 26144
rect 64396 26104 64436 26144
rect 64492 26104 64532 26144
rect 64684 26104 64724 26144
rect 64876 26104 64916 26144
rect 64972 26104 65012 26144
rect 65356 26104 65396 26144
rect 65548 26104 65588 26144
rect 65644 26104 65684 26144
rect 67180 26104 67220 26144
rect 67276 26104 67316 26144
rect 67372 26104 67412 26144
rect 67468 26104 67508 26144
rect 67660 26104 67700 26144
rect 67852 26104 67892 26144
rect 67948 26104 67988 26144
rect 68140 26104 68180 26144
rect 68332 26104 68372 26144
rect 69292 26104 69332 26144
rect 69388 26104 69428 26144
rect 69484 26104 69524 26144
rect 70924 26104 70964 26144
rect 71212 26104 71252 26144
rect 71788 26104 71828 26144
rect 71980 26104 72020 26144
rect 74188 26104 74228 26144
rect 74284 26104 74324 26144
rect 74476 26104 74516 26144
rect 74764 26104 74804 26144
rect 74860 26104 74900 26144
rect 74956 26104 74996 26144
rect 75148 26104 75188 26144
rect 75340 26104 75380 26144
rect 75436 26104 75476 26144
rect 76780 26104 76820 26144
rect 76972 26104 77012 26144
rect 77068 26104 77108 26144
rect 652 26020 692 26060
rect 36652 26020 36692 26060
rect 38860 26020 38900 26060
rect 40396 26020 40436 26060
rect 40972 26020 41012 26060
rect 51916 26020 51956 26060
rect 58828 26020 58868 26060
rect 60364 26020 60404 26060
rect 60556 26020 60596 26060
rect 60940 26020 60980 26060
rect 68812 26020 68852 26060
rect 70444 26020 70484 26060
rect 844 25936 884 25976
rect 31948 25936 31988 25976
rect 35308 25936 35348 25976
rect 36268 25936 36308 25976
rect 36844 25936 36884 25976
rect 37708 25936 37748 25976
rect 39724 25936 39764 25976
rect 42220 25936 42260 25976
rect 47404 25936 47444 25976
rect 52876 25936 52916 25976
rect 55084 25936 55124 25976
rect 55372 25936 55412 25976
rect 56812 25936 56852 25976
rect 57964 25936 58004 25976
rect 58348 25936 58388 25976
rect 60172 25936 60212 25976
rect 60748 25936 60788 25976
rect 65356 25936 65396 25976
rect 66412 25936 66452 25976
rect 68620 25936 68660 25976
rect 39244 25852 39284 25892
rect 40588 25852 40628 25892
rect 40780 25852 40820 25892
rect 46252 25852 46292 25892
rect 48364 25852 48404 25892
rect 51244 25852 51284 25892
rect 52108 25852 52148 25892
rect 52588 25852 52628 25892
rect 59020 25852 59060 25892
rect 59404 25852 59444 25892
rect 59980 25852 60020 25892
rect 64012 25852 64052 25892
rect 73420 25894 73460 25934
rect 74476 25936 74516 25976
rect 68236 25852 68276 25892
rect 71596 25852 71636 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 34732 25516 34772 25556
rect 35404 25516 35444 25556
rect 35692 25516 35732 25556
rect 40396 25516 40436 25556
rect 40876 25516 40916 25556
rect 44044 25516 44084 25556
rect 54796 25516 54836 25556
rect 67756 25516 67796 25556
rect 75628 25516 75668 25556
rect 30316 25432 30356 25472
rect 32716 25432 32756 25472
rect 41356 25432 41396 25472
rect 42796 25432 42836 25472
rect 43852 25432 43892 25472
rect 46348 25432 46388 25472
rect 51436 25432 51476 25472
rect 55564 25432 55604 25472
rect 63820 25432 63860 25472
rect 73036 25432 73076 25472
rect 75916 25432 75956 25472
rect 652 25348 692 25388
rect 40684 25348 40724 25388
rect 31948 25264 31988 25304
rect 32044 25264 32084 25304
rect 32140 25264 32180 25304
rect 33196 25264 33236 25304
rect 33388 25264 33428 25304
rect 33484 25264 33524 25304
rect 34252 25264 34292 25304
rect 34348 25264 34388 25304
rect 34444 25264 34484 25304
rect 34540 25264 34580 25304
rect 34732 25264 34772 25304
rect 34924 25264 34964 25304
rect 35020 25264 35060 25304
rect 35308 25264 35348 25304
rect 35500 25264 35540 25304
rect 35692 25264 35732 25304
rect 35884 25264 35924 25304
rect 35980 25264 36020 25304
rect 36364 25264 36404 25304
rect 37228 25264 37268 25304
rect 37612 25264 37652 25304
rect 38476 25264 38516 25304
rect 39820 25264 39860 25304
rect 39916 25264 39956 25304
rect 40012 25264 40052 25304
rect 40108 25264 40148 25304
rect 40300 25264 40340 25304
rect 40492 25264 40532 25304
rect 44044 25264 44084 25304
rect 44236 25264 44276 25304
rect 44332 25264 44372 25304
rect 44620 25264 44660 25304
rect 44716 25264 44756 25304
rect 44812 25264 44852 25304
rect 45964 25264 46004 25304
rect 46252 25264 46292 25304
rect 46444 25264 46484 25304
rect 46732 25264 46772 25304
rect 46924 25264 46964 25304
rect 47500 25264 47540 25304
rect 48364 25264 48404 25304
rect 50572 25264 50612 25304
rect 50668 25264 50708 25304
rect 50764 25264 50804 25304
rect 50860 25264 50900 25304
rect 51052 25264 51092 25304
rect 51244 25264 51284 25304
rect 51724 25264 51764 25304
rect 51820 25264 51860 25304
rect 52108 25264 52148 25304
rect 52780 25264 52820 25304
rect 53644 25264 53684 25304
rect 55756 25264 55796 25304
rect 55948 25264 55988 25304
rect 57484 25264 57524 25304
rect 57868 25264 57908 25304
rect 58732 25264 58772 25304
rect 60172 25264 60212 25304
rect 60556 25264 60596 25304
rect 61420 25264 61460 25304
rect 63148 25264 63188 25304
rect 63436 25264 63476 25304
rect 63532 25264 63572 25304
rect 64396 25264 64436 25304
rect 65260 25264 65300 25304
rect 67084 25264 67124 25304
rect 67372 25264 67412 25304
rect 67468 25264 67508 25304
rect 68332 25251 68372 25291
rect 69196 25264 69236 25304
rect 71020 25264 71060 25304
rect 71884 25264 71924 25304
rect 73228 25264 73268 25304
rect 73612 25264 73652 25304
rect 74476 25264 74516 25304
rect 75820 25264 75860 25304
rect 76012 25264 76052 25304
rect 76204 25264 76244 25304
rect 76396 25264 76436 25304
rect 76492 25264 76532 25304
rect 77068 25264 77108 25304
rect 77932 25264 77972 25304
rect 46828 25180 46868 25220
rect 47116 25180 47156 25220
rect 51148 25180 51188 25220
rect 52396 25180 52436 25220
rect 55852 25180 55892 25220
rect 64012 25180 64052 25220
rect 67948 25180 67988 25220
rect 70636 25180 70676 25220
rect 76300 25180 76340 25220
rect 76684 25180 76724 25220
rect 844 25096 884 25136
rect 32236 25096 32276 25136
rect 33292 25096 33332 25136
rect 39628 25096 39668 25136
rect 40876 25096 40916 25136
rect 44524 25096 44564 25136
rect 49516 25096 49556 25136
rect 54796 25096 54836 25136
rect 59884 25096 59924 25136
rect 62572 25096 62612 25136
rect 66412 25096 66452 25136
rect 70348 25096 70388 25136
rect 75628 25096 75668 25136
rect 79084 25096 79124 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 37516 24760 37556 24800
rect 45004 24760 45044 24800
rect 50188 24760 50228 24800
rect 58348 24760 58388 24800
rect 58924 24760 58964 24800
rect 60460 24760 60500 24800
rect 64012 24760 64052 24800
rect 67756 24760 67796 24800
rect 70828 24760 70868 24800
rect 74380 24760 74420 24800
rect 29836 24676 29876 24716
rect 32524 24676 32564 24716
rect 46444 24676 46484 24716
rect 30220 24592 30260 24632
rect 31084 24592 31124 24632
rect 32428 24592 32468 24632
rect 32620 24592 32660 24632
rect 32716 24592 32756 24632
rect 35116 24592 35156 24632
rect 35500 24592 35540 24632
rect 36364 24592 36404 24632
rect 39532 24592 39572 24632
rect 39820 24592 39860 24632
rect 39916 24592 39956 24632
rect 40396 24592 40436 24632
rect 40588 24592 40628 24632
rect 40684 24592 40724 24632
rect 40876 24592 40916 24632
rect 40972 24592 41012 24632
rect 41068 24592 41108 24632
rect 42316 24592 42356 24632
rect 42700 24592 42740 24632
rect 43564 24592 43604 24632
rect 44908 24592 44948 24632
rect 45100 24592 45140 24632
rect 45196 24592 45236 24632
rect 46540 24592 46580 24632
rect 46828 24592 46868 24632
rect 47116 24592 47156 24632
rect 50380 24634 50420 24674
rect 59404 24676 59444 24716
rect 60172 24676 60212 24716
rect 64492 24676 64532 24716
rect 68236 24676 68276 24716
rect 75820 24676 75860 24716
rect 76588 24676 76628 24716
rect 47308 24592 47348 24632
rect 47404 24592 47444 24632
rect 50572 24592 50612 24632
rect 50668 24592 50708 24632
rect 52108 24592 52148 24632
rect 52300 24592 52340 24632
rect 52396 24592 52436 24632
rect 55084 24592 55124 24632
rect 55468 24592 55508 24632
rect 56332 24592 56372 24632
rect 58060 24592 58100 24632
rect 58156 24592 58196 24632
rect 58252 24592 58292 24632
rect 59500 24592 59540 24632
rect 59788 24592 59828 24632
rect 60076 24592 60116 24632
rect 60268 24592 60308 24632
rect 63532 24592 63572 24632
rect 63628 24592 63668 24632
rect 63724 24592 63764 24632
rect 63916 24592 63956 24632
rect 64108 24592 64148 24632
rect 64204 24592 64244 24632
rect 64396 24592 64436 24632
rect 64588 24592 64628 24632
rect 67660 24592 67700 24632
rect 67852 24592 67892 24632
rect 67948 24592 67988 24632
rect 68140 24592 68180 24632
rect 68332 24592 68372 24632
rect 70732 24592 70772 24632
rect 70924 24592 70964 24632
rect 71020 24592 71060 24632
rect 71596 24592 71636 24632
rect 71692 24592 71732 24632
rect 71788 24592 71828 24632
rect 74284 24592 74324 24632
rect 74476 24592 74516 24632
rect 74572 24592 74612 24632
rect 75436 24592 75476 24632
rect 75724 24592 75764 24632
rect 76492 24592 76532 24632
rect 76684 24592 76724 24632
rect 652 24508 692 24548
rect 39052 24508 39092 24548
rect 49996 24508 50036 24548
rect 51340 24508 51380 24548
rect 57484 24508 57524 24548
rect 58732 24508 58772 24548
rect 60652 24508 60692 24548
rect 40204 24424 40244 24464
rect 46156 24424 46196 24464
rect 47116 24424 47156 24464
rect 47596 24424 47636 24464
rect 48460 24424 48500 24464
rect 51148 24424 51188 24464
rect 52108 24424 52148 24464
rect 52588 24424 52628 24464
rect 59116 24424 59156 24464
rect 60844 24424 60884 24464
rect 64780 24424 64820 24464
rect 68524 24424 68564 24464
rect 71212 24424 71252 24464
rect 76108 24424 76148 24464
rect 77164 24424 77204 24464
rect 844 24340 884 24380
rect 32236 24340 32276 24380
rect 39244 24340 39284 24380
rect 40396 24340 40436 24380
rect 44716 24340 44756 24380
rect 50188 24340 50228 24380
rect 50380 24340 50420 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 2188 24004 2228 24044
rect 35500 24004 35540 24044
rect 35884 24004 35924 24044
rect 43276 24004 43316 24044
rect 44428 24004 44468 24044
rect 55372 24004 55412 24044
rect 28684 23920 28724 23960
rect 32716 23920 32756 23960
rect 37036 23920 37076 23960
rect 45772 23920 45812 23960
rect 46924 23920 46964 23960
rect 652 23836 692 23876
rect 1804 23836 1844 23876
rect 1996 23836 2036 23876
rect 31468 23836 31508 23876
rect 30700 23752 30740 23792
rect 30892 23752 30932 23792
rect 30988 23752 31028 23792
rect 32044 23752 32084 23792
rect 32332 23752 32372 23792
rect 33484 23752 33524 23792
rect 34348 23752 34388 23792
rect 35884 23752 35924 23792
rect 36076 23752 36116 23792
rect 36172 23752 36212 23792
rect 36364 23752 36404 23792
rect 37324 23752 37364 23792
rect 38860 23752 38900 23792
rect 38956 23752 38996 23792
rect 39052 23752 39092 23792
rect 39340 23752 39380 23792
rect 39532 23752 39572 23792
rect 39628 23752 39668 23792
rect 40492 23752 40532 23792
rect 40684 23752 40724 23792
rect 41260 23752 41300 23792
rect 42124 23752 42164 23792
rect 43948 23752 43988 23792
rect 44044 23752 44084 23792
rect 44140 23752 44180 23792
rect 44236 23752 44276 23792
rect 44428 23752 44468 23792
rect 44620 23752 44660 23792
rect 44716 23752 44756 23792
rect 45100 23752 45140 23792
rect 45388 23752 45428 23792
rect 45484 23752 45524 23792
rect 45964 23752 46004 23792
rect 46060 23752 46100 23792
rect 46156 23752 46196 23792
rect 48364 23752 48404 23792
rect 49228 23752 49268 23792
rect 50572 23752 50612 23792
rect 50764 23752 50804 23792
rect 50860 23752 50900 23792
rect 51052 23752 51092 23792
rect 51244 23752 51284 23792
rect 51340 23752 51380 23792
rect 51724 23752 51764 23792
rect 52108 23752 52148 23792
rect 52972 23752 53012 23792
rect 54796 23752 54836 23792
rect 55084 23752 55124 23792
rect 55372 23752 55412 23792
rect 55564 23752 55604 23792
rect 55660 23752 55700 23792
rect 55852 23752 55892 23792
rect 56140 23752 56180 23792
rect 56428 23752 56468 23792
rect 56812 23752 56852 23792
rect 57292 23752 57332 23792
rect 57676 23752 57716 23792
rect 58060 23752 58100 23792
rect 58444 23752 58484 23792
rect 58924 23752 58964 23792
rect 59308 23752 59348 23792
rect 59692 23752 59732 23792
rect 60076 23752 60116 23792
rect 60460 23752 60500 23792
rect 60844 23752 60884 23792
rect 61324 23752 61364 23792
rect 61708 23752 61748 23792
rect 62092 23752 62132 23792
rect 62476 23752 62516 23792
rect 62860 23752 62900 23792
rect 63244 23752 63284 23792
rect 63724 23752 63764 23792
rect 64108 23752 64148 23792
rect 64492 23752 64532 23792
rect 64876 23752 64916 23792
rect 65260 23752 65300 23792
rect 65740 23752 65780 23792
rect 66124 23752 66164 23792
rect 66508 23752 66548 23792
rect 66892 23752 66932 23792
rect 67276 23752 67316 23792
rect 67756 23752 67796 23792
rect 68140 23752 68180 23792
rect 68524 23752 68564 23792
rect 68908 23752 68948 23792
rect 69292 23752 69332 23792
rect 69772 23752 69812 23792
rect 70156 23752 70196 23792
rect 70540 23752 70580 23792
rect 70924 23752 70964 23792
rect 71308 23752 71348 23792
rect 71692 23752 71732 23792
rect 72076 23752 72116 23792
rect 72460 23752 72500 23792
rect 72844 23752 72884 23792
rect 73324 23752 73364 23792
rect 73708 23752 73748 23792
rect 74092 23752 74132 23792
rect 74476 23752 74516 23792
rect 74860 23752 74900 23792
rect 75244 23752 75284 23792
rect 75628 23752 75668 23792
rect 76108 23752 76148 23792
rect 76972 23752 77012 23792
rect 77260 23752 77300 23792
rect 77452 23752 77492 23792
rect 77740 23752 77780 23792
rect 78124 23752 78164 23792
rect 78508 23752 78548 23792
rect 78796 23752 78836 23792
rect 79084 23752 79124 23792
rect 79372 23752 79412 23792
rect 32428 23668 32468 23708
rect 33100 23668 33140 23708
rect 40588 23668 40628 23708
rect 40876 23668 40916 23708
rect 47980 23668 48020 23708
rect 51148 23668 51188 23708
rect 844 23584 884 23624
rect 1612 23584 1652 23624
rect 30796 23584 30836 23624
rect 31660 23584 31700 23624
rect 39148 23584 39188 23624
rect 39436 23584 39476 23624
rect 43276 23584 43316 23624
rect 50380 23584 50420 23624
rect 50668 23584 50708 23624
rect 54124 23584 54164 23624
rect 54892 23584 54932 23624
rect 55180 23584 55220 23624
rect 55948 23584 55988 23624
rect 56236 23584 56276 23624
rect 56524 23584 56564 23624
rect 56908 23584 56948 23624
rect 57388 23584 57428 23624
rect 57772 23584 57812 23624
rect 58156 23584 58196 23624
rect 58540 23584 58580 23624
rect 59020 23584 59060 23624
rect 59404 23584 59444 23624
rect 59788 23584 59828 23624
rect 60172 23584 60212 23624
rect 60556 23584 60596 23624
rect 60940 23584 60980 23624
rect 61420 23584 61460 23624
rect 61804 23584 61844 23624
rect 62188 23584 62228 23624
rect 62572 23584 62612 23624
rect 62956 23584 62996 23624
rect 63340 23584 63380 23624
rect 63820 23584 63860 23624
rect 64204 23584 64244 23624
rect 64588 23584 64628 23624
rect 64972 23584 65012 23624
rect 65356 23584 65396 23624
rect 65836 23584 65876 23624
rect 66220 23584 66260 23624
rect 66604 23584 66644 23624
rect 66988 23584 67028 23624
rect 67372 23584 67412 23624
rect 67852 23584 67892 23624
rect 68236 23584 68276 23624
rect 68620 23584 68660 23624
rect 69004 23584 69044 23624
rect 69388 23584 69428 23624
rect 69868 23584 69908 23624
rect 70252 23584 70292 23624
rect 70636 23584 70676 23624
rect 71020 23584 71060 23624
rect 71404 23584 71444 23624
rect 71788 23584 71828 23624
rect 72172 23584 72212 23624
rect 72556 23584 72596 23624
rect 72940 23584 72980 23624
rect 73420 23584 73460 23624
rect 73804 23584 73844 23624
rect 74188 23584 74228 23624
rect 74572 23584 74612 23624
rect 74956 23584 74996 23624
rect 75340 23584 75380 23624
rect 75724 23584 75764 23624
rect 76204 23584 76244 23624
rect 76876 23584 76916 23624
rect 77164 23584 77204 23624
rect 77548 23584 77588 23624
rect 77836 23584 77876 23624
rect 78220 23584 78260 23624
rect 78604 23584 78644 23624
rect 78892 23584 78932 23624
rect 79180 23584 79220 23624
rect 79468 23584 79508 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 41068 23290 41108 23330
rect 31276 23248 31316 23288
rect 32812 23248 32852 23288
rect 35692 23248 35732 23288
rect 37900 23248 37940 23288
rect 40876 23248 40916 23288
rect 44716 23248 44756 23288
rect 48844 23248 48884 23288
rect 49516 23248 49556 23288
rect 49996 23248 50036 23288
rect 28204 23164 28244 23204
rect 32428 23164 32468 23204
rect 36652 23164 36692 23204
rect 37228 23164 37268 23204
rect 41356 23164 41396 23204
rect 50668 23164 50708 23204
rect 51244 23164 51284 23204
rect 51628 23164 51668 23204
rect 1516 23080 1556 23120
rect 1900 23080 1940 23120
rect 2092 23080 2132 23120
rect 28588 23080 28628 23120
rect 29452 23080 29492 23120
rect 31180 23080 31220 23120
rect 31372 23080 31412 23120
rect 31468 23080 31508 23120
rect 32332 23080 32372 23120
rect 32524 23080 32564 23120
rect 32716 23080 32756 23120
rect 32908 23080 32948 23120
rect 33004 23080 33044 23120
rect 33196 23080 33236 23120
rect 33292 23080 33332 23120
rect 33388 23080 33428 23120
rect 35788 23080 35828 23120
rect 35884 23080 35924 23120
rect 35980 23080 36020 23120
rect 36268 23080 36308 23120
rect 36556 23080 36596 23120
rect 37132 23080 37172 23120
rect 37324 23080 37364 23120
rect 37804 23080 37844 23120
rect 37996 23080 38036 23120
rect 38092 23080 38132 23120
rect 38476 23080 38516 23120
rect 38860 23080 38900 23120
rect 39724 23080 39764 23120
rect 41452 23080 41492 23120
rect 41740 23080 41780 23120
rect 44620 23080 44660 23120
rect 44812 23080 44852 23120
rect 44908 23080 44948 23120
rect 45484 23080 45524 23120
rect 45580 23080 45620 23120
rect 45676 23080 45716 23120
rect 45868 23080 45908 23120
rect 45964 23080 46004 23120
rect 46156 23069 46196 23109
rect 46444 23080 46484 23120
rect 46828 23080 46868 23120
rect 47692 23080 47732 23120
rect 49708 23080 49748 23120
rect 49804 23080 49844 23120
rect 49900 23080 49940 23120
rect 50284 23080 50324 23120
rect 50572 23080 50612 23120
rect 51148 23080 51188 23120
rect 51340 23080 51380 23120
rect 51532 23101 51572 23141
rect 51724 23080 51764 23120
rect 52588 23080 52628 23120
rect 52684 23080 52724 23120
rect 652 22996 692 23036
rect 42412 22996 42452 23036
rect 49324 22996 49364 23036
rect 1516 22912 1556 22952
rect 33580 22912 33620 22952
rect 35500 22912 35540 22952
rect 36940 22912 36980 22952
rect 42028 22912 42068 22952
rect 42796 22912 42836 22952
rect 50956 22912 50996 22952
rect 844 22828 884 22868
rect 1708 22828 1748 22868
rect 1900 22828 1940 22868
rect 30604 22828 30644 22868
rect 42604 22828 42644 22868
rect 46156 22828 46196 22868
rect 49516 22828 49556 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 34924 22492 34964 22532
rect 39052 22492 39092 22532
rect 43468 22492 43508 22532
rect 51244 22492 51284 22532
rect 52012 22492 52052 22532
rect 52396 22492 52436 22532
rect 52684 22492 52724 22532
rect 652 22408 692 22448
rect 31564 22408 31604 22448
rect 35596 22408 35636 22448
rect 38188 22408 38228 22448
rect 38860 22408 38900 22448
rect 40396 22408 40436 22448
rect 46444 22408 46484 22448
rect 48172 22408 48212 22448
rect 3244 22324 3284 22364
rect 28012 22324 28052 22364
rect 40204 22324 40244 22364
rect 49036 22324 49076 22364
rect 30316 22240 30356 22280
rect 30412 22240 30452 22280
rect 30508 22240 30548 22280
rect 30604 22240 30644 22280
rect 30892 22240 30932 22280
rect 31180 22240 31220 22280
rect 31276 22240 31316 22280
rect 31852 22240 31892 22280
rect 32044 22240 32084 22280
rect 32140 22240 32180 22280
rect 32908 22240 32948 22280
rect 33772 22240 33812 22280
rect 36172 22240 36212 22280
rect 37036 22240 37076 22280
rect 39052 22240 39092 22280
rect 39244 22240 39284 22280
rect 39340 22240 39380 22280
rect 40588 22240 40628 22280
rect 40780 22240 40820 22280
rect 40876 22240 40916 22280
rect 41452 22240 41492 22280
rect 42316 22240 42356 22280
rect 45100 22240 45140 22280
rect 45292 22240 45332 22280
rect 45388 22240 45428 22280
rect 45580 22240 45620 22280
rect 45772 22240 45812 22280
rect 48556 22240 48596 22280
rect 48652 22240 48692 22280
rect 48748 22240 48788 22280
rect 49420 22240 49460 22280
rect 49612 22240 49652 22280
rect 49708 22240 49748 22280
rect 50188 22240 50228 22280
rect 50380 22240 50420 22280
rect 51436 22240 51476 22280
rect 52108 22240 52148 22280
rect 52300 22240 52340 22280
rect 52588 22240 52628 22280
rect 32524 22156 32564 22196
rect 35788 22156 35828 22196
rect 41068 22156 41108 22196
rect 45676 22156 45716 22196
rect 50284 22156 50324 22196
rect 3436 22072 3476 22112
rect 28204 22072 28244 22112
rect 31948 22072 31988 22112
rect 34924 22072 34964 22112
rect 40684 22072 40724 22112
rect 45196 22072 45236 22112
rect 48844 22072 48884 22112
rect 49228 22072 49268 22112
rect 49516 22072 49556 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 3244 21736 3284 21776
rect 29452 21736 29492 21776
rect 36268 21736 36308 21776
rect 44716 21736 44756 21776
rect 31564 21652 31604 21692
rect 32140 21652 32180 21692
rect 41164 21652 41204 21692
rect 42316 21652 42356 21692
rect 51052 21652 51092 21692
rect 3052 21568 3092 21608
rect 3148 21568 3188 21608
rect 3340 21568 3380 21608
rect 27820 21568 27860 21608
rect 27916 21568 27956 21608
rect 28012 21568 28052 21608
rect 28108 21568 28148 21608
rect 28300 21568 28340 21608
rect 28492 21568 28532 21608
rect 28588 21568 28628 21608
rect 28876 21568 28916 21608
rect 29068 21568 29108 21608
rect 29356 21568 29396 21608
rect 29548 21568 29588 21608
rect 29644 21568 29684 21608
rect 31468 21568 31508 21608
rect 31660 21568 31700 21608
rect 32044 21568 32084 21608
rect 32236 21568 32276 21608
rect 36172 21568 36212 21608
rect 36364 21568 36404 21608
rect 36460 21568 36500 21608
rect 36652 21568 36692 21608
rect 36844 21568 36884 21608
rect 39052 21568 39092 21608
rect 39148 21568 39188 21608
rect 39244 21568 39284 21608
rect 39340 21568 39380 21608
rect 41068 21568 41108 21608
rect 41260 21568 41300 21608
rect 42700 21568 42740 21608
rect 43564 21568 43604 21608
rect 45004 21568 45044 21608
rect 45292 21568 45332 21608
rect 45388 21568 45428 21608
rect 45964 21568 46004 21608
rect 46348 21568 46388 21608
rect 47212 21568 47252 21608
rect 48844 21568 48884 21608
rect 49036 21568 49076 21608
rect 49132 21568 49172 21608
rect 49516 21568 49556 21608
rect 49612 21568 49652 21608
rect 49708 21568 49748 21608
rect 50188 21568 50228 21608
rect 50284 21568 50324 21608
rect 50572 21568 50612 21608
rect 50860 21568 50900 21608
rect 50956 21568 50996 21608
rect 51148 21568 51188 21608
rect 52588 21568 52628 21608
rect 52684 21568 52724 21608
rect 2860 21473 2900 21513
rect 3724 21484 3764 21524
rect 5740 21484 5780 21524
rect 5932 21484 5972 21524
rect 26860 21484 26900 21524
rect 27436 21484 27476 21524
rect 48364 21484 48404 21524
rect 5548 21400 5588 21440
rect 26476 21400 26516 21440
rect 27052 21400 27092 21440
rect 27628 21400 27668 21440
rect 29836 21400 29876 21440
rect 32812 21400 32852 21440
rect 33196 21400 33236 21440
rect 35788 21400 35828 21440
rect 36748 21400 36788 21440
rect 39532 21400 39572 21440
rect 49900 21400 49940 21440
rect 51340 21400 51380 21440
rect 2668 21316 2708 21356
rect 3532 21316 3572 21356
rect 6124 21316 6164 21356
rect 28300 21316 28340 21356
rect 28972 21316 29012 21356
rect 45676 21316 45716 21356
rect 48844 21316 48884 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 31660 20980 31700 21020
rect 46060 20980 46100 21020
rect 46348 20980 46388 21020
rect 50092 20980 50132 21020
rect 52684 20980 52724 21020
rect 652 20896 692 20936
rect 41740 20896 41780 20936
rect 32044 20812 32084 20852
rect 42892 20812 42932 20852
rect 43468 20812 43508 20852
rect 43660 20812 43700 20852
rect 44140 20812 44180 20852
rect 5452 20728 5492 20768
rect 26956 20728 26996 20768
rect 27820 20728 27860 20768
rect 28204 20728 28244 20768
rect 28684 20728 28724 20768
rect 28876 20728 28916 20768
rect 28972 20728 29012 20768
rect 29644 20728 29684 20768
rect 30508 20728 30548 20768
rect 32716 20728 32756 20768
rect 33580 20728 33620 20768
rect 35788 20728 35828 20768
rect 36652 20728 36692 20768
rect 38284 20728 38324 20768
rect 38380 20728 38420 20768
rect 38572 20728 38612 20768
rect 39148 20728 39188 20768
rect 40012 20728 40052 20768
rect 41932 20728 41972 20768
rect 42028 20728 42068 20768
rect 42220 20728 42260 20768
rect 44812 20728 44852 20768
rect 44908 20728 44948 20768
rect 45004 20728 45044 20768
rect 45100 20728 45140 20768
rect 45484 20728 45524 20768
rect 45676 20728 45716 20768
rect 45772 20728 45812 20768
rect 45964 20728 46004 20768
rect 46156 20728 46196 20768
rect 46348 20728 46388 20768
rect 46540 20728 46580 20768
rect 46636 20728 46676 20768
rect 47692 20728 47732 20768
rect 48076 20728 48116 20768
rect 48940 20728 48980 20768
rect 50284 20728 50324 20768
rect 50668 20728 50708 20768
rect 51532 20728 51572 20768
rect 28780 20644 28820 20684
rect 29260 20644 29300 20684
rect 32332 20644 32372 20684
rect 35404 20644 35444 20684
rect 38764 20644 38804 20684
rect 5548 20560 5588 20600
rect 25804 20560 25844 20600
rect 31852 20560 31892 20600
rect 34732 20560 34772 20600
rect 37804 20560 37844 20600
rect 38476 20560 38516 20600
rect 41164 20560 41204 20600
rect 42124 20560 42164 20600
rect 43084 20560 43124 20600
rect 43276 20560 43316 20600
rect 43852 20560 43892 20600
rect 44332 20560 44372 20600
rect 45580 20560 45620 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 35692 20224 35732 20264
rect 41164 20140 41204 20180
rect 41452 20140 41492 20180
rect 22732 20056 22772 20096
rect 22828 20056 22868 20096
rect 22924 20056 22964 20096
rect 23020 20056 23060 20096
rect 26668 20056 26708 20096
rect 26860 20056 26900 20096
rect 26956 20056 26996 20096
rect 27916 20056 27956 20096
rect 28204 20056 28244 20096
rect 28300 20056 28340 20096
rect 28780 20056 28820 20096
rect 28876 20056 28916 20096
rect 28983 20069 29023 20109
rect 31180 20056 31220 20096
rect 32044 20056 32084 20096
rect 32620 20056 32660 20096
rect 32716 20056 32756 20096
rect 32812 20056 32852 20096
rect 32908 20056 32948 20096
rect 33100 20041 33140 20081
rect 33292 20056 33332 20096
rect 34924 20056 34964 20096
rect 35020 20056 35060 20096
rect 35212 20056 35252 20096
rect 35500 20056 35540 20096
rect 35596 20056 35636 20096
rect 35788 20056 35828 20096
rect 35980 20056 36020 20096
rect 36076 20056 36116 20096
rect 36172 20056 36212 20096
rect 36268 20056 36308 20096
rect 37516 20056 37556 20096
rect 37708 20056 37748 20096
rect 37900 20056 37940 20096
rect 37996 20056 38036 20096
rect 38188 20056 38228 20096
rect 38572 20056 38612 20096
rect 40972 20056 41012 20096
rect 41068 20056 41108 20096
rect 41260 20056 41300 20096
rect 41836 20056 41876 20096
rect 42700 20056 42740 20096
rect 9004 19972 9044 20012
rect 22348 19972 22388 20012
rect 25612 19972 25652 20012
rect 26284 19972 26324 20012
rect 27148 19972 27188 20012
rect 44332 19972 44372 20012
rect 45292 19972 45332 20012
rect 45676 19972 45716 20012
rect 47500 19972 47540 20012
rect 47884 19972 47924 20012
rect 49324 19972 49364 20012
rect 652 19888 692 19928
rect 23308 19888 23348 19928
rect 26476 19888 26516 19928
rect 27340 19888 27380 19928
rect 28588 19888 28628 19928
rect 29740 19888 29780 19928
rect 35212 19888 35252 19928
rect 38188 19888 38228 19928
rect 44524 19888 44564 19928
rect 44716 19888 44756 19928
rect 46828 19888 46868 19928
rect 50092 19888 50132 19928
rect 9196 19804 9236 19844
rect 22540 19804 22580 19844
rect 25420 19804 25460 19844
rect 26668 19804 26708 19844
rect 31660 19804 31700 19844
rect 33196 19804 33236 19844
rect 37612 19804 37652 19844
rect 40108 19804 40148 19844
rect 43852 19804 43892 19844
rect 45100 19804 45140 19844
rect 45484 19804 45524 19844
rect 47308 19804 47348 19844
rect 47692 19804 47732 19844
rect 49132 19804 49172 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 11692 19468 11732 19508
rect 22156 19468 22196 19508
rect 32428 19468 32468 19508
rect 32908 19468 32948 19508
rect 35788 19468 35828 19508
rect 39052 19468 39092 19508
rect 652 19384 692 19424
rect 6604 19384 6644 19424
rect 8812 19384 8852 19424
rect 25900 19384 25940 19424
rect 33868 19384 33908 19424
rect 36076 19384 36116 19424
rect 38284 19384 38324 19424
rect 40300 19384 40340 19424
rect 40684 19384 40724 19424
rect 43564 19384 43604 19424
rect 21580 19300 21620 19340
rect 21964 19300 22004 19340
rect 37228 19300 37268 19340
rect 41260 19300 41300 19340
rect 41644 19300 41684 19340
rect 42028 19300 42068 19340
rect 8332 19216 8372 19256
rect 8524 19216 8564 19256
rect 8620 19216 8660 19256
rect 8812 19216 8852 19256
rect 9004 19216 9044 19256
rect 9100 19216 9140 19256
rect 9292 19216 9332 19256
rect 9676 19216 9716 19256
rect 10540 19216 10580 19256
rect 22348 19216 22388 19256
rect 22444 19216 22484 19256
rect 22636 19202 22676 19242
rect 23212 19216 23252 19256
rect 24076 19216 24116 19256
rect 26476 19216 26516 19256
rect 27373 19216 27413 19256
rect 29644 19216 29684 19256
rect 30508 19216 30548 19256
rect 32140 19216 32180 19256
rect 32236 19216 32276 19256
rect 32428 19216 32468 19256
rect 33196 19216 33236 19256
rect 33292 19216 33332 19256
rect 33580 19216 33620 19256
rect 35692 19216 35732 19256
rect 35884 19216 35924 19256
rect 36364 19216 36404 19256
rect 36460 19216 36500 19256
rect 36748 19216 36788 19256
rect 38188 19216 38228 19256
rect 38380 19216 38420 19256
rect 38572 19216 38612 19256
rect 38668 19216 38708 19256
rect 38860 19216 38900 19256
rect 39340 19216 39380 19256
rect 39436 19216 39476 19256
rect 39724 19216 39764 19256
rect 42220 19216 42260 19256
rect 42316 19216 42356 19256
rect 42412 19216 42452 19256
rect 42508 19216 42548 19256
rect 42892 19216 42932 19256
rect 43180 19189 43220 19229
rect 43276 19216 43316 19256
rect 44140 19216 44180 19256
rect 45004 19216 45044 19256
rect 46732 19216 46772 19256
rect 47596 19216 47636 19256
rect 49036 19216 49076 19256
rect 49228 19216 49268 19256
rect 49324 19216 49364 19256
rect 49996 19216 50036 19256
rect 50860 19216 50900 19256
rect 22828 19132 22868 19172
rect 26092 19132 26132 19172
rect 29260 19132 29300 19172
rect 43756 19132 43796 19172
rect 46348 19132 46388 19172
rect 49132 19132 49172 19172
rect 49612 19132 49652 19172
rect 8428 19048 8468 19088
rect 11692 19048 11732 19088
rect 21772 19048 21812 19088
rect 22156 19048 22196 19088
rect 22540 19048 22580 19088
rect 25228 19048 25268 19088
rect 28492 19048 28532 19088
rect 31660 19048 31700 19088
rect 37036 19048 37076 19088
rect 38764 19048 38804 19088
rect 41068 19048 41108 19088
rect 41452 19048 41492 19088
rect 41836 19048 41876 19088
rect 46156 19048 46196 19088
rect 48748 19048 48788 19088
rect 52012 19048 52052 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 9004 18712 9044 18752
rect 26092 18712 26132 18752
rect 29356 18712 29396 18752
rect 42892 18712 42932 18752
rect 44044 18712 44084 18752
rect 8332 18628 8372 18668
rect 8812 18628 8852 18668
rect 9484 18628 9524 18668
rect 23116 18628 23156 18668
rect 30604 18628 30644 18668
rect 32620 18628 32660 18668
rect 35788 18628 35828 18668
rect 36172 18628 36212 18668
rect 38764 18628 38804 18668
rect 48076 18628 48116 18668
rect 48652 18628 48692 18668
rect 49420 18628 49460 18668
rect 7084 18544 7124 18584
rect 7948 18544 7988 18584
rect 8524 18544 8564 18584
rect 8716 18544 8756 18584
rect 8620 18502 8660 18542
rect 9388 18544 9428 18584
rect 9580 18544 9620 18584
rect 22732 18544 22772 18584
rect 23020 18544 23060 18584
rect 25324 18544 25364 18584
rect 25420 18544 25460 18584
rect 25612 18544 25652 18584
rect 25900 18544 25940 18584
rect 25996 18544 26036 18584
rect 26188 18544 26228 18584
rect 26380 18544 26420 18584
rect 26476 18544 26516 18584
rect 26572 18544 26612 18584
rect 26668 18544 26708 18584
rect 28684 18544 28724 18584
rect 28780 18544 28820 18584
rect 28972 18544 29012 18584
rect 29164 18544 29204 18584
rect 29260 18544 29300 18584
rect 29452 18544 29492 18584
rect 29644 18544 29684 18584
rect 29740 18544 29780 18584
rect 29836 18544 29876 18584
rect 29932 18544 29972 18584
rect 30220 18544 30260 18584
rect 30508 18544 30548 18584
rect 31084 18544 31124 18584
rect 31276 18544 31316 18584
rect 31852 18544 31892 18584
rect 31948 18544 31988 18584
rect 32140 18544 32180 18584
rect 32524 18544 32564 18584
rect 32716 18544 32756 18584
rect 32812 18544 32852 18584
rect 33004 18544 33044 18584
rect 33388 18544 33428 18584
rect 34252 18544 34292 18584
rect 35692 18544 35732 18584
rect 35884 18544 35924 18584
rect 35980 18544 36020 18584
rect 36556 18544 36596 18584
rect 37420 18544 37460 18584
rect 39148 18544 39188 18584
rect 39964 18544 40004 18584
rect 41932 18544 41972 18584
rect 42124 18544 42164 18584
rect 42220 18544 42260 18584
rect 42412 18544 42452 18584
rect 42604 18544 42644 18584
rect 42700 18544 42740 18584
rect 43564 18544 43604 18584
rect 43660 18544 43700 18584
rect 43756 18544 43796 18584
rect 43948 18544 43988 18584
rect 44140 18544 44180 18584
rect 44236 18544 44276 18584
rect 44428 18544 44468 18584
rect 44524 18544 44564 18584
rect 44620 18544 44660 18584
rect 46156 18544 46196 18584
rect 46348 18544 46388 18584
rect 46732 18544 46772 18584
rect 46828 18544 46868 18584
rect 47020 18544 47060 18584
rect 47404 18544 47444 18584
rect 47500 18544 47540 18584
rect 47596 18544 47636 18584
rect 47692 18544 47732 18584
rect 47980 18544 48020 18584
rect 48172 18544 48212 18584
rect 48748 18544 48788 18584
rect 49036 18544 49076 18584
rect 49324 18544 49364 18584
rect 49516 18544 49556 18584
rect 52300 18544 52340 18584
rect 52684 18544 52724 18584
rect 9196 18460 9236 18500
rect 21484 18460 21524 18500
rect 22060 18460 22100 18500
rect 22252 18460 22292 18500
rect 23596 18460 23636 18500
rect 23980 18460 24020 18500
rect 24364 18460 24404 18500
rect 41164 18460 41204 18500
rect 41740 18460 41780 18500
rect 43084 18460 43124 18500
rect 49900 18460 49940 18500
rect 50572 18460 50612 18500
rect 51340 18460 51380 18500
rect 652 18376 692 18416
rect 9772 18376 9812 18416
rect 23788 18376 23828 18416
rect 25612 18376 25652 18416
rect 28972 18376 29012 18416
rect 30892 18376 30932 18416
rect 32140 18376 32180 18416
rect 42412 18376 42452 18416
rect 46252 18376 46292 18416
rect 48364 18376 48404 18416
rect 50764 18376 50804 18416
rect 5932 18292 5972 18332
rect 9004 18292 9044 18332
rect 21676 18292 21716 18332
rect 21868 18292 21908 18332
rect 22444 18292 22484 18332
rect 23404 18292 23444 18332
rect 24172 18292 24212 18332
rect 24556 18292 24596 18332
rect 31180 18292 31220 18332
rect 35404 18292 35444 18332
rect 38572 18292 38612 18332
rect 41548 18292 41588 18332
rect 41932 18292 41972 18332
rect 42892 18292 42932 18332
rect 47020 18292 47060 18332
rect 50092 18292 50132 18332
rect 50380 18292 50420 18332
rect 51148 18292 51188 18332
rect 52396 18292 52436 18332
rect 52588 18292 52628 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 8620 17956 8660 17996
rect 22444 17956 22484 17996
rect 26476 17956 26516 17996
rect 33388 17956 33428 17996
rect 36460 17956 36500 17996
rect 46348 17956 46388 17996
rect 652 17872 692 17912
rect 8332 17872 8372 17912
rect 26764 17872 26804 17912
rect 27724 17872 27764 17912
rect 34732 17872 34772 17912
rect 36748 17872 36788 17912
rect 37804 17872 37844 17912
rect 48460 17872 48500 17912
rect 50092 17872 50132 17912
rect 1708 17788 1748 17828
rect 22252 17788 22292 17828
rect 46540 17788 46580 17828
rect 48268 17788 48308 17828
rect 49420 17788 49460 17828
rect 7660 17704 7700 17744
rect 7948 17704 7988 17744
rect 8524 17704 8564 17744
rect 8716 17704 8756 17744
rect 22636 17704 22676 17744
rect 22828 17704 22868 17744
rect 22924 17704 22964 17744
rect 23500 17704 23540 17744
rect 24364 17704 24404 17744
rect 26380 17704 26420 17744
rect 26572 17704 26612 17744
rect 27052 17704 27092 17744
rect 27148 17704 27188 17744
rect 27436 17704 27476 17744
rect 29932 17704 29972 17744
rect 30124 17704 30164 17744
rect 30220 17704 30260 17744
rect 30796 17704 30836 17744
rect 31660 17704 31700 17744
rect 33292 17704 33332 17744
rect 33484 17704 33524 17744
rect 34156 17704 34196 17744
rect 34348 17704 34388 17744
rect 36364 17704 36404 17744
rect 36556 17704 36596 17744
rect 39820 17704 39860 17744
rect 40204 17704 40244 17744
rect 41068 17704 41108 17744
rect 42700 17704 42740 17744
rect 42892 17704 42932 17744
rect 42988 17704 43028 17744
rect 43564 17704 43604 17744
rect 44428 17704 44468 17744
rect 46060 17704 46100 17744
rect 46156 17704 46196 17744
rect 46348 17704 46388 17744
rect 48652 17704 48692 17744
rect 48748 17704 48788 17744
rect 48940 17704 48980 17744
rect 49804 17704 49844 17744
rect 49900 17718 49940 17758
rect 50092 17704 50132 17744
rect 50284 17704 50324 17744
rect 50668 17704 50708 17744
rect 51532 17704 51572 17744
rect 8044 17620 8084 17660
rect 22732 17620 22772 17660
rect 23116 17620 23156 17660
rect 30028 17620 30068 17660
rect 30412 17620 30452 17660
rect 34252 17620 34292 17660
rect 42796 17620 42836 17660
rect 43180 17620 43220 17660
rect 1516 17536 1556 17576
rect 25516 17536 25556 17576
rect 32812 17536 32852 17576
rect 42220 17536 42260 17576
rect 45580 17536 45620 17576
rect 46732 17536 46772 17576
rect 48844 17536 48884 17576
rect 49612 17536 49652 17576
rect 52684 17536 52724 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 2476 17200 2516 17240
rect 26860 17200 26900 17240
rect 41644 17200 41684 17240
rect 22828 17116 22868 17156
rect 23212 17116 23252 17156
rect 27244 17116 27284 17156
rect 33868 17116 33908 17156
rect 44140 17116 44180 17156
rect 45772 17116 45812 17156
rect 51340 17116 51380 17156
rect 22732 17032 22772 17072
rect 22924 17032 22964 17072
rect 23116 17032 23156 17072
rect 23308 17032 23348 17072
rect 26764 17032 26804 17072
rect 26956 17032 26996 17072
rect 27052 17032 27092 17072
rect 27628 17032 27668 17072
rect 28492 17032 28532 17072
rect 30508 17032 30548 17072
rect 30700 17032 30740 17072
rect 33772 17032 33812 17072
rect 33964 17032 34004 17072
rect 34060 17032 34100 17072
rect 34252 17032 34292 17072
rect 34636 17032 34676 17072
rect 35500 17032 35540 17072
rect 36940 17032 36980 17072
rect 37132 17032 37172 17072
rect 37324 17032 37364 17072
rect 37708 17032 37748 17072
rect 38572 17032 38612 17072
rect 41740 17032 41780 17072
rect 41836 17032 41876 17072
rect 41932 17032 41972 17072
rect 42220 17032 42260 17072
rect 42508 17032 42548 17072
rect 42604 17032 42644 17072
rect 44044 17032 44084 17072
rect 44236 17032 44276 17072
rect 45388 17032 45428 17072
rect 45676 17032 45716 17072
rect 46252 17032 46292 17072
rect 46636 17032 46676 17072
rect 47500 17032 47540 17072
rect 49132 17032 49172 17072
rect 49228 17032 49268 17072
rect 49420 17032 49460 17072
rect 50380 17032 50420 17072
rect 50668 17032 50708 17072
rect 50764 17032 50804 17072
rect 51244 17032 51284 17072
rect 51436 17032 51476 17072
rect 52300 17032 52340 17072
rect 52588 17032 52628 17072
rect 2668 16948 2708 16988
rect 33388 16948 33428 16988
rect 41068 16948 41108 16988
rect 41452 16948 41492 16988
rect 43084 16948 43124 16988
rect 44524 16948 44564 16988
rect 44908 16948 44948 16988
rect 48652 16948 48692 16988
rect 49900 16948 49940 16988
rect 51628 16961 51668 17001
rect 52396 16948 52436 16988
rect 652 16864 692 16904
rect 23692 16864 23732 16904
rect 30604 16864 30644 16904
rect 30892 16864 30932 16904
rect 36652 16864 36692 16904
rect 40876 16864 40916 16904
rect 42892 16864 42932 16904
rect 43660 16864 43700 16904
rect 44716 16864 44756 16904
rect 52684 16864 52724 16904
rect 29644 16780 29684 16820
rect 33580 16780 33620 16820
rect 37036 16780 37076 16820
rect 39724 16780 39764 16820
rect 41260 16780 41300 16820
rect 43276 16780 43316 16820
rect 45100 16780 45140 16820
rect 46060 16780 46100 16820
rect 49420 16780 49460 16820
rect 50092 16780 50132 16820
rect 51052 16780 51092 16820
rect 51820 16780 51860 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 4204 16444 4244 16484
rect 34636 16444 34676 16484
rect 37996 16444 38036 16484
rect 42700 16444 42740 16484
rect 42988 16444 43028 16484
rect 45676 16444 45716 16484
rect 45964 16444 46004 16484
rect 51340 16444 51380 16484
rect 54508 16444 54548 16484
rect 54892 16444 54932 16484
rect 55756 16444 55796 16484
rect 56236 16444 56276 16484
rect 56620 16444 56660 16484
rect 57388 16444 57428 16484
rect 58060 16444 58100 16484
rect 58348 16444 58388 16484
rect 58636 16444 58676 16484
rect 60172 16444 60212 16484
rect 60652 16444 60692 16484
rect 61516 16444 61556 16484
rect 62188 16444 62228 16484
rect 62476 16444 62516 16484
rect 63052 16444 63092 16484
rect 63340 16444 63380 16484
rect 63628 16444 63668 16484
rect 63916 16444 63956 16484
rect 64588 16444 64628 16484
rect 65068 16444 65108 16484
rect 65452 16444 65492 16484
rect 65836 16444 65876 16484
rect 66604 16444 66644 16484
rect 67084 16444 67124 16484
rect 67468 16444 67508 16484
rect 67852 16444 67892 16484
rect 68236 16444 68276 16484
rect 69100 16444 69140 16484
rect 69484 16444 69524 16484
rect 69868 16444 69908 16484
rect 70252 16444 70292 16484
rect 70636 16444 70676 16484
rect 71020 16444 71060 16484
rect 71404 16444 71444 16484
rect 71884 16444 71924 16484
rect 72268 16444 72308 16484
rect 72652 16444 72692 16484
rect 73036 16444 73076 16484
rect 73420 16444 73460 16484
rect 74284 16444 74324 16484
rect 74668 16444 74708 16484
rect 75052 16444 75092 16484
rect 75436 16444 75476 16484
rect 75820 16444 75860 16484
rect 76492 16444 76532 16484
rect 76876 16444 76916 16484
rect 77260 16444 77300 16484
rect 77548 16444 77588 16484
rect 77932 16444 77972 16484
rect 78316 16444 78356 16484
rect 78700 16444 78740 16484
rect 78988 16444 79028 16484
rect 79276 16444 79316 16484
rect 652 16360 692 16400
rect 1516 16360 1556 16400
rect 2380 16360 2420 16400
rect 34348 16360 34388 16400
rect 36748 16360 36788 16400
rect 46828 16360 46868 16400
rect 53164 16360 53204 16400
rect 53644 16360 53684 16400
rect 57580 16360 57620 16400
rect 61036 16360 61076 16400
rect 1996 16276 2036 16316
rect 2572 16276 2612 16316
rect 2764 16276 2804 16316
rect 4396 16276 4436 16316
rect 46636 16276 46676 16316
rect 61708 16276 61748 16316
rect 3340 16192 3380 16232
rect 3532 16192 3572 16232
rect 4972 16192 5012 16232
rect 5836 16192 5876 16232
rect 27353 16207 27393 16247
rect 27532 16192 27572 16232
rect 31372 16192 31412 16232
rect 32236 16192 32276 16232
rect 33676 16192 33716 16232
rect 33964 16192 34004 16232
rect 34540 16192 34580 16232
rect 34732 16192 34772 16232
rect 36364 16192 36404 16232
rect 36460 16192 36500 16232
rect 36556 16192 36596 16232
rect 37132 16192 37172 16232
rect 37420 16192 37460 16232
rect 37708 16192 37748 16232
rect 37804 16192 37844 16232
rect 37996 16192 38036 16232
rect 39916 16192 39956 16232
rect 40108 16192 40148 16232
rect 40684 16192 40724 16232
rect 41548 16192 41588 16232
rect 42892 16192 42932 16232
rect 43084 16192 43124 16232
rect 43660 16192 43700 16232
rect 44524 16192 44564 16232
rect 45964 16192 46004 16232
rect 46156 16192 46196 16232
rect 46252 16192 46292 16232
rect 48652 16192 48692 16232
rect 49036 16192 49076 16232
rect 49900 16192 49940 16232
rect 51244 16192 51284 16232
rect 51436 16192 51476 16232
rect 51628 16192 51668 16232
rect 52588 16192 52628 16232
rect 52780 16192 52820 16232
rect 52876 16192 52916 16232
rect 53068 16192 53108 16232
rect 53269 16179 53309 16219
rect 54412 16192 54452 16232
rect 54796 16192 54836 16232
rect 55276 16192 55316 16232
rect 55660 16192 55700 16232
rect 56140 16192 56180 16232
rect 56524 16192 56564 16232
rect 56908 16192 56948 16232
rect 57292 16192 57332 16232
rect 57964 16192 58004 16232
rect 58252 16192 58292 16232
rect 58540 16192 58580 16232
rect 58924 16192 58964 16232
rect 59308 16192 59348 16232
rect 59692 16192 59732 16232
rect 60076 16192 60116 16232
rect 60556 16192 60596 16232
rect 61420 16192 61460 16232
rect 62092 16192 62132 16232
rect 62380 16192 62420 16232
rect 62668 16192 62708 16232
rect 62956 16192 62996 16232
rect 63244 16192 63284 16232
rect 63532 16192 63572 16232
rect 63820 16192 63860 16232
rect 64108 16192 64148 16232
rect 64492 16192 64532 16232
rect 64972 16192 65012 16232
rect 65356 16192 65396 16232
rect 65740 16192 65780 16232
rect 66124 16192 66164 16232
rect 66508 16192 66548 16232
rect 66988 16192 67028 16232
rect 67372 16192 67412 16232
rect 67756 16192 67796 16232
rect 68140 16192 68180 16232
rect 68524 16192 68564 16232
rect 69004 16192 69044 16232
rect 69388 16192 69428 16232
rect 69772 16192 69812 16232
rect 70156 16192 70196 16232
rect 70527 16181 70567 16221
rect 70924 16192 70964 16232
rect 71308 16192 71348 16232
rect 71788 16192 71828 16232
rect 72172 16192 72212 16232
rect 72556 16192 72596 16232
rect 72940 16192 72980 16232
rect 73324 16192 73364 16232
rect 73708 16192 73748 16232
rect 74188 16192 74228 16232
rect 74572 16192 74612 16232
rect 74956 16192 74996 16232
rect 75340 16192 75380 16232
rect 75724 16192 75764 16232
rect 76588 16192 76628 16232
rect 76972 16192 77012 16232
rect 77164 16192 77204 16232
rect 77452 16192 77492 16232
rect 77836 16192 77876 16232
rect 78220 16192 78260 16232
rect 78604 16192 78644 16232
rect 78892 16192 78932 16232
rect 79180 16192 79220 16232
rect 3436 16108 3476 16148
rect 4588 16108 4628 16148
rect 27436 16108 27476 16148
rect 30988 16108 31028 16148
rect 34060 16108 34100 16148
rect 37036 16108 37076 16148
rect 40012 16108 40052 16148
rect 40300 16108 40340 16148
rect 43276 16108 43316 16148
rect 55372 16108 55412 16148
rect 2188 16024 2228 16064
rect 2956 16024 2996 16064
rect 6988 16024 7028 16064
rect 33388 16024 33428 16064
rect 45676 16024 45716 16064
rect 46444 16024 46484 16064
rect 51052 16024 51092 16064
rect 52684 16024 52724 16064
rect 57004 16024 57044 16064
rect 59020 16024 59060 16064
rect 59404 16024 59444 16064
rect 59788 16024 59828 16064
rect 61900 16024 61940 16064
rect 62764 16024 62804 16064
rect 64204 16024 64244 16064
rect 66220 16024 66260 16064
rect 68620 16024 68660 16064
rect 73804 16024 73844 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 3628 15688 3668 15728
rect 4396 15688 4436 15728
rect 33868 15688 33908 15728
rect 34924 15688 34964 15728
rect 40492 15688 40532 15728
rect 45964 15688 46004 15728
rect 49708 15688 49748 15728
rect 59500 15688 59540 15728
rect 67852 15688 67892 15728
rect 70540 15688 70580 15728
rect 79468 15688 79508 15728
rect 53164 15604 53204 15644
rect 1036 15520 1076 15560
rect 1420 15520 1460 15560
rect 2284 15520 2324 15560
rect 4204 15520 4244 15560
rect 4300 15520 4340 15560
rect 4492 15520 4532 15560
rect 4684 15520 4724 15560
rect 4780 15520 4820 15560
rect 4876 15520 4916 15560
rect 31948 15520 31988 15560
rect 32140 15520 32180 15560
rect 32812 15520 32852 15560
rect 33004 15520 33044 15560
rect 33118 15520 33158 15560
rect 33292 15520 33332 15560
rect 33388 15520 33428 15560
rect 33484 15520 33524 15560
rect 33580 15520 33620 15560
rect 33772 15520 33812 15560
rect 33964 15520 34004 15560
rect 34060 15520 34100 15560
rect 34444 15520 34484 15560
rect 34636 15520 34676 15560
rect 34732 15520 34772 15560
rect 36076 15520 36116 15560
rect 36940 15520 36980 15560
rect 37324 15520 37364 15560
rect 37516 15520 37556 15560
rect 37708 15520 37748 15560
rect 37804 15520 37844 15560
rect 39052 15520 39092 15560
rect 39148 15520 39188 15560
rect 39244 15520 39284 15560
rect 39724 15520 39764 15560
rect 39820 15520 39860 15560
rect 40108 15520 40148 15560
rect 40396 15520 40436 15560
rect 40588 15520 40628 15560
rect 40684 15520 40724 15560
rect 41836 15520 41876 15560
rect 42028 15520 42068 15560
rect 42124 15520 42164 15560
rect 45388 15520 45428 15560
rect 45484 15520 45524 15560
rect 45580 15520 45620 15560
rect 45676 15520 45716 15560
rect 45868 15520 45908 15560
rect 46060 15520 46100 15560
rect 46156 15520 46196 15560
rect 46348 15520 46388 15560
rect 46444 15520 46484 15560
rect 46540 15520 46580 15560
rect 46924 15520 46964 15560
rect 47212 15478 47252 15518
rect 47308 15520 47348 15560
rect 47788 15520 47828 15560
rect 47980 15520 48020 15560
rect 49804 15520 49844 15560
rect 49900 15520 49940 15560
rect 49996 15520 50036 15560
rect 50850 15527 50890 15567
rect 50956 15520 50996 15560
rect 51148 15520 51188 15560
rect 51532 15520 51572 15560
rect 51628 15520 51668 15560
rect 51724 15520 51764 15560
rect 51820 15520 51860 15560
rect 52204 15520 52244 15560
rect 52492 15520 52532 15560
rect 52588 15520 52628 15560
rect 53548 15520 53588 15560
rect 54412 15520 54452 15560
rect 57100 15520 57140 15560
rect 57484 15520 57524 15560
rect 58348 15520 58388 15560
rect 60556 15520 60596 15560
rect 60940 15520 60980 15560
rect 61804 15520 61844 15560
rect 64780 15520 64820 15560
rect 64972 15520 65012 15560
rect 65452 15520 65492 15560
rect 65836 15520 65876 15560
rect 66700 15520 66740 15560
rect 70060 15520 70100 15560
rect 70156 15520 70196 15560
rect 70348 15520 70388 15560
rect 75148 15520 75188 15560
rect 75340 15520 75380 15560
rect 79372 15520 79412 15560
rect 844 15436 884 15476
rect 3820 15436 3860 15476
rect 55564 15436 55604 15476
rect 68716 15436 68756 15476
rect 69868 15436 69908 15476
rect 70732 15436 70772 15476
rect 71116 15436 71156 15476
rect 5068 15352 5108 15392
rect 31468 15352 31508 15392
rect 34444 15352 34484 15392
rect 37516 15352 37556 15392
rect 38188 15352 38228 15392
rect 39436 15352 39476 15392
rect 40876 15352 40916 15392
rect 43756 15352 43796 15392
rect 48460 15352 48500 15392
rect 49132 15352 49172 15392
rect 68044 15352 68084 15392
rect 71308 15352 71348 15392
rect 72652 15352 72692 15392
rect 76684 15352 76724 15392
rect 652 15268 692 15308
rect 3436 15268 3476 15308
rect 3628 15268 3668 15308
rect 32044 15268 32084 15308
rect 32812 15268 32852 15308
rect 41836 15268 41876 15308
rect 47596 15268 47636 15308
rect 47884 15268 47924 15308
rect 51148 15268 51188 15308
rect 52876 15268 52916 15308
rect 59500 15268 59540 15308
rect 62956 15268 62996 15308
rect 64876 15268 64916 15308
rect 68908 15268 68948 15308
rect 69676 15268 69716 15308
rect 70348 15268 70388 15308
rect 70924 15268 70964 15308
rect 75244 15268 75284 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 1996 14932 2036 14972
rect 3244 14932 3284 14972
rect 45580 14932 45620 14972
rect 50380 14932 50420 14972
rect 53164 14932 53204 14972
rect 56908 14932 56948 14972
rect 60940 14932 60980 14972
rect 65356 14932 65396 14972
rect 72748 14932 72788 14972
rect 75340 14932 75380 14972
rect 78604 14932 78644 14972
rect 652 14848 692 14888
rect 33484 14848 33524 14888
rect 35596 14848 35636 14888
rect 40012 14848 40052 14888
rect 45100 14848 45140 14888
rect 54316 14848 54356 14888
rect 56716 14848 56756 14888
rect 57484 14848 57524 14888
rect 58636 14848 58676 14888
rect 61420 14848 61460 14888
rect 64108 14848 64148 14888
rect 65932 14848 65972 14888
rect 844 14764 884 14804
rect 1228 14764 1268 14804
rect 60748 14764 60788 14804
rect 61612 14764 61652 14804
rect 61996 14764 62036 14804
rect 62764 14764 62804 14804
rect 67180 14764 67220 14804
rect 1516 14680 1556 14720
rect 1612 14680 1652 14720
rect 1708 14680 1748 14720
rect 1804 14680 1844 14720
rect 1996 14680 2036 14720
rect 2860 14722 2900 14762
rect 2188 14680 2228 14720
rect 2284 14680 2324 14720
rect 2572 14680 2612 14720
rect 2956 14680 2996 14720
rect 5068 14680 5108 14720
rect 5260 14680 5300 14720
rect 30316 14680 30356 14720
rect 31180 14680 31220 14720
rect 32812 14680 32852 14720
rect 32908 14680 32948 14720
rect 33004 14659 33044 14699
rect 35980 14680 36020 14720
rect 36076 14680 36116 14720
rect 36172 14680 36212 14720
rect 36268 14680 36308 14720
rect 36844 14680 36884 14720
rect 38572 14680 38612 14720
rect 39436 14680 39476 14720
rect 39820 14680 39860 14720
rect 40012 14680 40052 14720
rect 40204 14680 40244 14720
rect 40300 14680 40340 14720
rect 41260 14680 41300 14720
rect 41356 14680 41396 14720
rect 41452 14680 41492 14720
rect 42796 14680 42836 14720
rect 42988 14680 43028 14720
rect 43084 14680 43124 14720
rect 43276 14680 43316 14720
rect 43372 14680 43412 14720
rect 43468 14680 43508 14720
rect 45580 14680 45620 14720
rect 45772 14680 45812 14720
rect 45868 14680 45908 14720
rect 46252 14680 46292 14720
rect 47404 14680 47444 14720
rect 47596 14680 47636 14720
rect 48364 14680 48404 14720
rect 49228 14680 49268 14720
rect 51148 14680 51188 14720
rect 52012 14680 52052 14720
rect 56044 14680 56084 14720
rect 56332 14680 56372 14720
rect 56908 14680 56948 14720
rect 57100 14680 57140 14720
rect 57196 14680 57236 14720
rect 57388 14680 57428 14720
rect 57580 14680 57620 14720
rect 60940 14680 60980 14720
rect 61132 14680 61172 14720
rect 61228 14680 61268 14720
rect 62188 14680 62228 14720
rect 62284 14680 62324 14720
rect 62380 14680 62420 14720
rect 63724 14680 63764 14720
rect 63820 14680 63860 14720
rect 63916 14680 63956 14720
rect 64492 14680 64532 14720
rect 64780 14680 64820 14720
rect 65068 14680 65108 14720
rect 65164 14680 65204 14720
rect 65356 14680 65396 14720
rect 67948 14680 67988 14720
rect 68812 14680 68852 14720
rect 70348 14680 70388 14720
rect 70732 14680 70772 14720
rect 71596 14680 71636 14720
rect 73612 14680 73652 14720
rect 73804 14680 73844 14720
rect 73900 14680 73940 14720
rect 74092 14680 74132 14720
rect 74188 14680 74228 14720
rect 74284 14680 74324 14720
rect 74380 14680 74420 14720
rect 74668 14680 74708 14720
rect 74956 14680 74996 14720
rect 75628 14680 75668 14720
rect 75820 14680 75860 14720
rect 75916 14680 75956 14720
rect 76204 14680 76244 14720
rect 76588 14680 76628 14720
rect 77452 14680 77492 14720
rect 5164 14596 5204 14636
rect 29932 14596 29972 14636
rect 47500 14596 47540 14636
rect 47980 14596 48020 14636
rect 50764 14596 50804 14636
rect 56428 14596 56468 14636
rect 64396 14596 64436 14636
rect 67564 14596 67604 14636
rect 75052 14596 75092 14636
rect 75724 14596 75764 14636
rect 1036 14512 1076 14552
rect 32332 14512 32372 14552
rect 32716 14512 32756 14552
rect 37420 14512 37460 14552
rect 41548 14512 41588 14552
rect 42892 14512 42932 14552
rect 53164 14512 53204 14552
rect 60556 14512 60596 14552
rect 61804 14512 61844 14552
rect 62572 14512 62612 14552
rect 67372 14512 67412 14552
rect 69964 14512 70004 14552
rect 72748 14512 72788 14552
rect 73708 14512 73748 14552
rect 78604 14512 78644 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 1132 14176 1172 14216
rect 2380 14176 2420 14216
rect 2860 14176 2900 14216
rect 7468 14176 7508 14216
rect 35404 14176 35444 14216
rect 38380 14176 38420 14216
rect 39436 14176 39476 14216
rect 51340 14176 51380 14216
rect 52108 14176 52148 14216
rect 56236 14176 56276 14216
rect 68524 14176 68564 14216
rect 69004 14176 69044 14216
rect 70540 14176 70580 14216
rect 79372 14176 79412 14216
rect 32332 14092 32372 14132
rect 40012 14092 40052 14132
rect 43180 14092 43220 14132
rect 47692 14092 47732 14132
rect 52972 14092 53012 14132
rect 68236 14092 68276 14132
rect 2764 14008 2804 14048
rect 2956 14008 2996 14048
rect 3052 14008 3092 14048
rect 4012 14008 4052 14048
rect 4300 14008 4340 14048
rect 4396 14008 4436 14048
rect 5068 14008 5108 14048
rect 5452 14008 5492 14048
rect 6316 14008 6356 14048
rect 31468 14008 31508 14048
rect 31660 14008 31700 14048
rect 31756 14008 31796 14048
rect 32428 14008 32468 14048
rect 32716 14008 32756 14048
rect 33004 14008 33044 14048
rect 33388 14008 33428 14048
rect 34252 14008 34292 14048
rect 37228 14008 37268 14048
rect 38092 14008 38132 14048
rect 38284 14008 38324 14048
rect 38476 14008 38516 14048
rect 38572 14008 38612 14048
rect 39148 14008 39188 14048
rect 39244 14008 39284 14048
rect 39340 14008 39380 14048
rect 39820 14008 39860 14048
rect 39916 14008 39956 14048
rect 40108 14008 40148 14048
rect 40300 14008 40340 14048
rect 40684 14008 40724 14048
rect 41548 14008 41588 14048
rect 43276 14008 43316 14048
rect 43564 14008 43604 14048
rect 44620 14008 44660 14048
rect 45004 14008 45044 14048
rect 45868 14008 45908 14048
rect 47596 14008 47636 14048
rect 47788 14008 47828 14048
rect 47884 14008 47924 14048
rect 51148 14008 51188 14048
rect 51244 14008 51284 14048
rect 51436 14008 51476 14048
rect 52588 14008 52628 14048
rect 52876 14008 52916 14048
rect 53068 14008 53108 14048
rect 53356 14008 53396 14048
rect 53452 14008 53492 14048
rect 53644 14008 53684 14048
rect 53836 14008 53876 14048
rect 54220 14008 54260 14048
rect 55084 14008 55124 14048
rect 56428 14008 56468 14048
rect 56620 14008 56660 14048
rect 57772 14008 57812 14048
rect 57964 14008 58004 14048
rect 58156 14008 58196 14048
rect 58540 14008 58580 14048
rect 59404 14008 59444 14048
rect 60844 14008 60884 14048
rect 61036 14008 61076 14048
rect 61228 14008 61268 14048
rect 61612 14008 61652 14048
rect 62476 14008 62516 14048
rect 63820 14008 63860 14048
rect 63916 14008 63956 14048
rect 64108 14008 64148 14048
rect 64684 14008 64724 14048
rect 65068 14008 65108 14048
rect 65932 14008 65972 14048
rect 67276 14008 67316 14048
rect 67372 14008 67412 14048
rect 67564 14008 67604 14048
rect 68044 14008 68084 14048
rect 68140 14008 68180 14048
rect 68332 14050 68372 14090
rect 70060 14092 70100 14132
rect 71020 14092 71060 14132
rect 72172 14092 72212 14132
rect 75916 14092 75956 14132
rect 68620 14029 68660 14069
rect 68716 14008 68756 14048
rect 68812 14008 68852 14048
rect 69676 14008 69716 14048
rect 69964 14008 70004 14048
rect 70924 14008 70964 14048
rect 71116 14008 71156 14048
rect 72556 14008 72596 14048
rect 73420 13997 73460 14037
rect 74764 14008 74804 14048
rect 74956 14008 74996 14048
rect 75052 14008 75092 14048
rect 75820 14008 75860 14048
rect 76012 14008 76052 14048
rect 76972 14008 77012 14048
rect 77356 14008 77396 14048
rect 78220 14008 78260 14048
rect 1324 13924 1364 13964
rect 1708 13924 1748 13964
rect 2572 13924 2612 13964
rect 47020 13924 47060 13964
rect 67084 13924 67124 13964
rect 69196 13924 69236 13964
rect 70732 13924 70772 13964
rect 30412 13840 30452 13880
rect 31468 13840 31508 13880
rect 43852 13840 43892 13880
rect 50956 13840 50996 13880
rect 67564 13840 67604 13880
rect 1516 13756 1556 13796
rect 4684 13756 4724 13796
rect 32044 13756 32084 13796
rect 37612 13756 37652 13796
rect 42700 13756 42740 13796
rect 42892 13756 42932 13796
rect 53644 13756 53684 13796
rect 56236 13756 56276 13796
rect 56524 13756 56564 13796
rect 57868 13756 57908 13796
rect 60556 13756 60596 13796
rect 60940 13756 60980 13796
rect 63628 13756 63668 13796
rect 64108 13756 64148 13796
rect 70348 13756 70388 13796
rect 74572 13756 74612 13796
rect 74764 13756 74804 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 4492 13420 4532 13460
rect 32428 13420 32468 13460
rect 33004 13420 33044 13460
rect 36268 13420 36308 13460
rect 41548 13420 41588 13460
rect 42796 13420 42836 13460
rect 45484 13420 45524 13460
rect 47308 13420 47348 13460
rect 54700 13420 54740 13460
rect 58732 13420 58772 13460
rect 61036 13420 61076 13460
rect 64588 13420 64628 13460
rect 70156 13420 70196 13460
rect 76492 13420 76532 13460
rect 1228 13336 1268 13376
rect 1900 13336 1940 13376
rect 5356 13336 5396 13376
rect 6220 13336 6260 13376
rect 39532 13336 39572 13376
rect 40780 13336 40820 13376
rect 51820 13336 51860 13376
rect 56332 13336 56372 13376
rect 58540 13336 58580 13376
rect 62476 13336 62516 13376
rect 65164 13336 65204 13376
rect 71020 13336 71060 13376
rect 71980 13336 72020 13376
rect 74572 13336 74612 13376
rect 76108 13336 76148 13376
rect 77068 13336 77108 13376
rect 77452 13336 77492 13376
rect 844 13252 884 13292
rect 1420 13252 1460 13292
rect 6700 13252 6740 13292
rect 1612 13168 1652 13208
rect 1708 13168 1748 13208
rect 1900 13168 1940 13208
rect 2092 13168 2132 13208
rect 2476 13168 2516 13208
rect 3340 13168 3380 13208
rect 5164 13168 5204 13208
rect 6028 13168 6068 13208
rect 6604 13168 6644 13208
rect 6796 13168 6836 13208
rect 32332 13168 32372 13208
rect 32524 13168 32564 13208
rect 32716 13168 32756 13208
rect 32812 13168 32852 13208
rect 33004 13168 33044 13208
rect 34828 13168 34868 13208
rect 34924 13168 34964 13208
rect 35116 13168 35156 13208
rect 36172 13191 36212 13231
rect 36364 13168 36404 13208
rect 36556 13168 36596 13208
rect 36748 13168 36788 13208
rect 37324 13168 37364 13208
rect 38188 13168 38228 13208
rect 41548 13168 41588 13208
rect 41740 13168 41780 13208
rect 41836 13168 41876 13208
rect 42700 13168 42740 13208
rect 42892 13168 42932 13208
rect 43084 13168 43124 13208
rect 43468 13168 43508 13208
rect 44332 13168 44372 13208
rect 46156 13168 46196 13208
rect 47308 13168 47348 13208
rect 47500 13182 47540 13222
rect 47596 13168 47636 13208
rect 47884 13168 47924 13208
rect 48076 13210 48116 13250
rect 47980 13168 48020 13208
rect 48652 13168 48692 13208
rect 48844 13168 48884 13208
rect 49804 13168 49844 13208
rect 50668 13168 50708 13208
rect 54412 13168 54452 13208
rect 54508 13168 54548 13208
rect 54700 13168 54740 13208
rect 55084 13168 55124 13208
rect 55180 13168 55220 13208
rect 55276 13168 55316 13208
rect 55372 13168 55412 13208
rect 56044 13168 56084 13208
rect 56140 13168 56180 13208
rect 56332 13168 56372 13208
rect 56524 13168 56564 13208
rect 56716 13168 56756 13208
rect 56812 13168 56852 13208
rect 57868 13168 57908 13208
rect 58156 13168 58196 13208
rect 58732 13168 58772 13208
rect 58924 13168 58964 13208
rect 59020 13168 59060 13208
rect 61324 13168 61364 13208
rect 61420 13168 61460 13208
rect 61708 13168 61748 13208
rect 62092 13168 62132 13208
rect 62188 13168 62228 13208
rect 62284 13168 62324 13208
rect 63916 13168 63956 13208
rect 64012 13168 64052 13208
rect 64108 13168 64148 13208
rect 64300 13168 64340 13208
rect 64396 13168 64436 13208
rect 64588 13168 64628 13208
rect 68716 13168 68756 13208
rect 68812 13168 68852 13208
rect 68908 13168 68948 13208
rect 69100 13168 69140 13208
rect 69292 13168 69332 13208
rect 69388 13168 69428 13208
rect 69676 13168 69716 13208
rect 69868 13168 69908 13208
rect 70060 13168 70100 13208
rect 70252 13168 70292 13208
rect 72172 13168 72212 13208
rect 72556 13168 72596 13208
rect 73420 13179 73460 13219
rect 74764 13168 74804 13208
rect 74860 13168 74900 13208
rect 74956 13168 74996 13208
rect 75052 13168 75092 13208
rect 75436 13168 75476 13208
rect 75724 13168 75764 13208
rect 75820 13168 75860 13208
rect 76492 13168 76532 13208
rect 76684 13168 76724 13208
rect 76780 13168 76820 13208
rect 76972 13168 77012 13208
rect 77164 13168 77204 13208
rect 36652 13084 36692 13124
rect 36940 13084 36980 13124
rect 48748 13084 48788 13124
rect 49420 13084 49460 13124
rect 58252 13084 58292 13124
rect 69772 13084 69812 13124
rect 652 13000 692 13040
rect 35020 13000 35060 13040
rect 39340 13000 39380 13040
rect 46636 13000 46676 13040
rect 48172 13000 48212 13040
rect 56620 13000 56660 13040
rect 61996 13000 62036 13040
rect 63820 13000 63860 13040
rect 68620 13000 68660 13040
rect 69196 13000 69236 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 1900 12664 1940 12704
rect 4588 12664 4628 12704
rect 41452 12664 41492 12704
rect 47884 12664 47924 12704
rect 49132 12664 49172 12704
rect 57292 12664 57332 12704
rect 61420 12664 61460 12704
rect 67180 12664 67220 12704
rect 72844 12664 72884 12704
rect 74380 12664 74420 12704
rect 48556 12580 48596 12620
rect 54892 12580 54932 12620
rect 1996 12517 2036 12557
rect 2092 12517 2132 12557
rect 844 12412 884 12452
rect 1324 12412 1364 12452
rect 1708 12412 1748 12452
rect 2188 12451 2228 12491
rect 2380 12496 2420 12536
rect 2572 12496 2612 12536
rect 2668 12496 2708 12536
rect 4492 12496 4532 12536
rect 4684 12496 4724 12536
rect 4780 12496 4820 12536
rect 5356 12496 5396 12536
rect 33868 12496 33908 12536
rect 34252 12496 34292 12536
rect 35116 12496 35156 12536
rect 36748 12496 36788 12536
rect 36844 12496 36884 12536
rect 37132 12496 37172 12536
rect 39052 12496 39092 12536
rect 39436 12496 39476 12536
rect 40300 12496 40340 12536
rect 42220 12496 42260 12536
rect 42412 12496 42452 12536
rect 45484 12496 45524 12536
rect 45868 12496 45908 12536
rect 46732 12496 46772 12536
rect 48172 12496 48212 12536
rect 48460 12496 48500 12536
rect 49036 12496 49076 12536
rect 49228 12496 49268 12536
rect 49324 12496 49364 12536
rect 49516 12496 49556 12536
rect 49612 12496 49652 12536
rect 49708 12496 49748 12536
rect 51628 12496 51668 12536
rect 51820 12496 51860 12536
rect 52012 12496 52052 12536
rect 52396 12496 52436 12536
rect 53260 12496 53300 12536
rect 55276 12496 55316 12536
rect 56140 12496 56180 12536
rect 58252 12496 58292 12536
rect 58444 12496 58484 12536
rect 59308 12496 59348 12536
rect 59500 12496 59540 12536
rect 61324 12496 61364 12536
rect 61516 12496 61556 12536
rect 61612 12496 61652 12536
rect 62092 12496 62132 12536
rect 62284 12496 62324 12536
rect 62380 12496 62420 12536
rect 63052 12496 63092 12536
rect 63244 12496 63284 12536
rect 63340 12496 63380 12536
rect 64396 12496 64436 12536
rect 64588 12496 64628 12536
rect 64780 12496 64820 12536
rect 65164 12496 65204 12536
rect 66028 12496 66068 12536
rect 67372 12496 67412 12536
rect 67756 12496 67796 12536
rect 68620 12496 68660 12536
rect 69964 12496 70004 12536
rect 70060 12496 70100 12536
rect 70252 12496 70292 12536
rect 70444 12496 70484 12536
rect 70828 12496 70868 12536
rect 71692 12496 71732 12536
rect 74284 12496 74324 12536
rect 74764 12538 74804 12578
rect 76108 12580 76148 12620
rect 74476 12496 74516 12536
rect 74572 12496 74612 12536
rect 74956 12496 74996 12536
rect 75052 12496 75092 12536
rect 76012 12496 76052 12536
rect 76204 12496 76244 12536
rect 76876 12496 76916 12536
rect 77260 12496 77300 12536
rect 78124 12496 78164 12536
rect 36268 12412 36308 12452
rect 54412 12412 54452 12452
rect 57868 12412 57908 12452
rect 652 12328 692 12368
rect 1132 12328 1172 12368
rect 2380 12328 2420 12368
rect 2860 12328 2900 12368
rect 5932 12328 5972 12368
rect 36460 12328 36500 12368
rect 37420 12328 37460 12368
rect 42796 12328 42836 12368
rect 48844 12328 48884 12368
rect 49900 12328 49940 12368
rect 58348 12328 58388 12368
rect 59788 12328 59828 12368
rect 62092 12328 62132 12368
rect 70252 12328 70292 12368
rect 74764 12328 74804 12368
rect 1516 12244 1556 12284
rect 42316 12244 42356 12284
rect 51724 12244 51764 12284
rect 58060 12244 58100 12284
rect 59404 12244 59444 12284
rect 63052 12244 63092 12284
rect 64492 12244 64532 12284
rect 69772 12244 69812 12284
rect 79276 12244 79316 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 34828 11908 34868 11948
rect 36844 11908 36884 11948
rect 39436 11908 39476 11948
rect 44716 11908 44756 11948
rect 46828 11908 46868 11948
rect 48268 11908 48308 11948
rect 61708 11908 61748 11948
rect 64588 11908 64628 11948
rect 69484 11908 69524 11948
rect 70540 11908 70580 11948
rect 74860 11908 74900 11948
rect 76396 11908 76436 11948
rect 1228 11824 1268 11864
rect 1804 11824 1844 11864
rect 4012 11824 4052 11864
rect 34348 11824 34388 11864
rect 38476 11824 38516 11864
rect 42124 11824 42164 11864
rect 44908 11824 44948 11864
rect 45964 11824 46004 11864
rect 49132 11824 49172 11864
rect 49804 11824 49844 11864
rect 51436 11824 51476 11864
rect 52492 11824 52532 11864
rect 55372 11824 55412 11864
rect 56332 11824 56372 11864
rect 57292 11824 57332 11864
rect 62092 11824 62132 11864
rect 64108 11824 64148 11864
rect 65356 11824 65396 11864
rect 67564 11824 67604 11864
rect 76012 11824 76052 11864
rect 77356 11824 77396 11864
rect 844 11740 884 11780
rect 1420 11740 1460 11780
rect 7372 11740 7412 11780
rect 49612 11740 49652 11780
rect 57484 11740 57524 11780
rect 1996 11656 2036 11696
rect 2092 11656 2132 11696
rect 2188 11656 2228 11696
rect 3340 11656 3380 11696
rect 3628 11656 3668 11696
rect 3724 11656 3764 11696
rect 4492 11656 4532 11696
rect 4684 11656 4724 11696
rect 4780 11656 4820 11696
rect 4972 11656 5012 11696
rect 5356 11656 5396 11696
rect 6220 11656 6260 11696
rect 34828 11656 34868 11696
rect 35020 11656 35060 11696
rect 35116 11656 35156 11696
rect 35308 11656 35348 11696
rect 35404 11656 35444 11696
rect 35500 11656 35540 11696
rect 35596 11656 35636 11696
rect 36076 11656 36116 11696
rect 36172 11656 36212 11696
rect 36364 11656 36404 11696
rect 36556 11656 36596 11696
rect 36652 11656 36692 11696
rect 36844 11656 36884 11696
rect 38092 11656 38132 11696
rect 38284 11656 38324 11696
rect 38860 11656 38900 11696
rect 39148 11656 39188 11696
rect 39436 11656 39476 11696
rect 39628 11656 39668 11696
rect 39724 11656 39764 11696
rect 41836 11656 41876 11696
rect 41932 11656 41972 11696
rect 42124 11656 42164 11696
rect 42316 11656 42356 11696
rect 42700 11656 42740 11696
rect 43564 11656 43604 11696
rect 46348 11656 46388 11696
rect 46444 11656 46484 11696
rect 46540 11656 46580 11696
rect 46636 11656 46676 11696
rect 46828 11656 46868 11696
rect 47020 11656 47060 11696
rect 47116 11656 47156 11696
rect 48268 11656 48308 11696
rect 48460 11656 48500 11696
rect 48556 11656 48596 11696
rect 49132 11656 49172 11696
rect 49324 11656 49364 11696
rect 49420 11656 49460 11696
rect 50188 11635 50228 11675
rect 50284 11656 50324 11696
rect 50380 11656 50420 11696
rect 50764 11656 50804 11696
rect 51052 11656 51092 11696
rect 51628 11656 51668 11696
rect 51724 11656 51764 11696
rect 51916 11656 51956 11696
rect 53740 11656 53780 11696
rect 53932 11656 53972 11696
rect 56524 11656 56564 11696
rect 56620 11656 56660 11696
rect 56716 11656 56756 11696
rect 56812 11656 56852 11696
rect 57676 11656 57716 11696
rect 57868 11656 57908 11696
rect 57964 11656 58004 11696
rect 58252 11656 58292 11696
rect 58348 11656 58388 11696
rect 58444 11656 58484 11696
rect 58828 11656 58868 11696
rect 59020 11656 59060 11696
rect 59116 11656 59156 11696
rect 59692 11656 59732 11696
rect 60556 11656 60596 11696
rect 62764 11635 62804 11675
rect 62860 11656 62900 11696
rect 62956 11656 62996 11696
rect 63052 11656 63092 11696
rect 63436 11656 63476 11696
rect 63724 11656 63764 11696
rect 64300 11656 64340 11696
rect 64396 11656 64436 11696
rect 64588 11656 64628 11696
rect 68908 11656 68948 11696
rect 69100 11656 69140 11696
rect 69196 11656 69236 11696
rect 69868 11656 69908 11696
rect 70156 11656 70196 11696
rect 70444 11656 70484 11696
rect 70636 11656 70676 11696
rect 72844 11656 72884 11696
rect 73708 11656 73748 11696
rect 75340 11656 75380 11696
rect 75628 11656 75668 11696
rect 75724 11656 75764 11696
rect 76396 11656 76436 11696
rect 76588 11656 76628 11696
rect 76684 11656 76724 11696
rect 76876 11656 76916 11696
rect 77068 11656 77108 11696
rect 4588 11572 4628 11612
rect 38188 11572 38228 11612
rect 38764 11572 38804 11612
rect 51148 11572 51188 11612
rect 51820 11572 51860 11612
rect 53836 11572 53876 11612
rect 58924 11572 58964 11612
rect 59308 11572 59348 11612
rect 63820 11572 63860 11612
rect 69004 11572 69044 11612
rect 69772 11572 69812 11612
rect 72460 11572 72500 11612
rect 76972 11572 77012 11612
rect 652 11488 692 11528
rect 2284 11488 2324 11528
rect 36268 11488 36308 11528
rect 50476 11488 50516 11528
rect 57772 11488 57812 11528
rect 58156 11488 58196 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 3916 11152 3956 11192
rect 37804 11152 37844 11192
rect 50476 11152 50516 11192
rect 56236 11152 56276 11192
rect 58828 11152 58868 11192
rect 60940 11152 60980 11192
rect 75244 11152 75284 11192
rect 4972 11068 5012 11108
rect 47020 11068 47060 11108
rect 48076 11068 48116 11108
rect 50860 11068 50900 11108
rect 59308 11068 59348 11108
rect 63340 11068 63380 11108
rect 64012 11068 64052 11108
rect 76204 11068 76244 11108
rect 1516 10984 1556 11024
rect 1900 10984 1940 11024
rect 2764 10984 2804 11024
rect 4108 10984 4148 11024
rect 4300 10984 4340 11024
rect 4876 10984 4916 11024
rect 5068 10984 5108 11024
rect 36364 10984 36404 11024
rect 36460 10984 36500 11024
rect 36652 10984 36692 11024
rect 36844 10984 36884 11024
rect 36940 10984 36980 11024
rect 37036 10984 37076 11024
rect 37132 10984 37172 11024
rect 39436 10984 39476 11024
rect 41548 10984 41588 11024
rect 41836 10984 41876 11024
rect 41932 10984 41972 11024
rect 42412 10984 42452 11024
rect 42604 10984 42644 11024
rect 43276 10984 43316 11024
rect 43468 10984 43508 11024
rect 43660 10984 43700 11024
rect 43756 10984 43796 11024
rect 43948 10984 43988 11024
rect 44140 10984 44180 11024
rect 44524 10984 44564 11024
rect 45388 10984 45428 11024
rect 46924 10984 46964 11024
rect 47116 10984 47156 11024
rect 48460 10984 48500 11024
rect 49324 10984 49364 11024
rect 50764 10984 50804 11024
rect 50956 10984 50996 11024
rect 51052 10984 51092 11024
rect 51340 10984 51380 11024
rect 51532 10984 51572 11024
rect 53356 10984 53396 11024
rect 53548 10984 53588 11024
rect 53644 10984 53684 11024
rect 53836 10984 53876 11024
rect 54220 10984 54260 11024
rect 55084 10984 55124 11024
rect 56428 10984 56468 11024
rect 56812 10984 56852 11024
rect 57676 10984 57716 11024
rect 59404 10984 59444 11024
rect 59692 10984 59732 11024
rect 62092 10984 62132 11024
rect 62956 10984 62996 11024
rect 63916 10984 63956 11024
rect 64108 10984 64148 11024
rect 64588 10984 64628 11024
rect 64780 10984 64820 11024
rect 64972 10984 65012 11024
rect 65164 10984 65204 11024
rect 65260 10984 65300 11024
rect 69004 10984 69044 11024
rect 69196 10984 69236 11024
rect 69292 10984 69332 11024
rect 74668 10984 74708 11024
rect 74764 10984 74804 11024
rect 74860 10984 74900 11024
rect 74956 10984 74996 11024
rect 75148 10984 75188 11024
rect 75340 10984 75380 11024
rect 75436 10984 75476 11024
rect 75628 10984 75668 11024
rect 75820 10984 75860 11024
rect 75916 10984 75956 11024
rect 76108 10984 76148 11024
rect 76300 10984 76340 11024
rect 77059 10997 77099 11037
rect 77260 10984 77300 11024
rect 844 10900 884 10940
rect 1324 10900 1364 10940
rect 51916 10900 51956 10940
rect 68812 10900 68852 10940
rect 69676 10900 69716 10940
rect 70156 10900 70196 10940
rect 70540 10900 70580 10940
rect 71116 10900 71156 10940
rect 76492 10900 76532 10940
rect 1132 10816 1172 10856
rect 36172 10816 36212 10856
rect 39820 10816 39860 10856
rect 42220 10816 42260 10856
rect 43372 10816 43412 10856
rect 43948 10816 43988 10856
rect 46540 10816 46580 10856
rect 47884 10816 47924 10856
rect 51436 10816 51476 10856
rect 65836 10816 65876 10856
rect 71308 10816 71348 10856
rect 72940 10816 72980 10856
rect 75628 10816 75668 10856
rect 77644 10816 77684 10856
rect 652 10732 692 10772
rect 4204 10732 4244 10772
rect 36652 10732 36692 10772
rect 42508 10732 42548 10772
rect 51724 10732 51764 10772
rect 53356 10732 53396 10772
rect 59020 10732 59060 10772
rect 64684 10732 64724 10772
rect 64972 10732 65012 10772
rect 68620 10732 68660 10772
rect 69004 10732 69044 10772
rect 69484 10732 69524 10772
rect 69964 10732 70004 10772
rect 70732 10732 70772 10772
rect 70924 10732 70964 10772
rect 76684 10732 76724 10772
rect 77164 10732 77204 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 38764 10396 38804 10436
rect 41740 10396 41780 10436
rect 49132 10396 49172 10436
rect 58060 10396 58100 10436
rect 63436 10396 63476 10436
rect 64972 10396 65012 10436
rect 67660 10396 67700 10436
rect 72844 10396 72884 10436
rect 75820 10396 75860 10436
rect 76876 10396 76916 10436
rect 1516 10312 1556 10352
rect 2188 10312 2228 10352
rect 2668 10312 2708 10352
rect 3148 10312 3188 10352
rect 5260 10312 5300 10352
rect 44140 10312 44180 10352
rect 53356 10312 53396 10352
rect 54316 10312 54356 10352
rect 57580 10312 57620 10352
rect 58732 10312 58772 10352
rect 60268 10312 60308 10352
rect 62380 10312 62420 10352
rect 67852 10312 67892 10352
rect 69964 10312 70004 10352
rect 844 10228 884 10268
rect 1708 10228 1748 10268
rect 3340 10228 3380 10268
rect 42124 10228 42164 10268
rect 57388 10228 57428 10268
rect 58924 10228 58964 10268
rect 59500 10228 59540 10268
rect 60076 10228 60116 10268
rect 79468 10228 79508 10268
rect 2188 10144 2228 10184
rect 2380 10144 2420 10184
rect 2476 10144 2516 10184
rect 2668 10144 2708 10184
rect 2956 10144 2996 10184
rect 36364 10144 36404 10184
rect 2860 10102 2900 10142
rect 36748 10144 36788 10184
rect 37612 10144 37652 10184
rect 38956 10144 38996 10184
rect 39148 10144 39188 10184
rect 39724 10144 39764 10184
rect 40588 10144 40628 10184
rect 43468 10144 43508 10184
rect 43756 10144 43796 10184
rect 44332 10144 44372 10184
rect 44524 10144 44564 10184
rect 46252 10144 46292 10184
rect 46444 10144 46484 10184
rect 46540 10144 46580 10184
rect 47116 10144 47156 10184
rect 47980 10144 48020 10184
rect 50284 10144 50324 10184
rect 51148 10144 51188 10184
rect 52684 10144 52724 10184
rect 52972 10144 53012 10184
rect 53548 10144 53588 10184
rect 53740 10144 53780 10184
rect 57772 10144 57812 10184
rect 57868 10144 57908 10184
rect 58060 10144 58100 10184
rect 58252 10144 58292 10184
rect 58444 10144 58484 10184
rect 58540 10144 58580 10184
rect 59116 10144 59156 10184
rect 59308 10144 59348 10184
rect 63436 10144 63476 10184
rect 63628 10144 63668 10184
rect 63724 10144 63764 10184
rect 64300 10144 64340 10184
rect 64588 10144 64628 10184
rect 65260 10144 65300 10184
rect 65644 10144 65684 10184
rect 66508 10144 66548 10184
rect 68236 10144 68276 10184
rect 68332 10144 68372 10184
rect 68428 10144 68468 10184
rect 68524 10144 68564 10184
rect 68716 10144 68756 10184
rect 68908 10144 68948 10184
rect 69004 10144 69044 10184
rect 69292 10144 69332 10184
rect 69580 10144 69620 10184
rect 69676 10144 69716 10184
rect 70828 10144 70868 10184
rect 71692 10144 71732 10184
rect 73804 10144 73844 10184
rect 74668 10144 74708 10184
rect 76204 10144 76244 10184
rect 76492 10144 76532 10184
rect 76588 10144 76628 10184
rect 77452 10144 77492 10184
rect 78316 10144 78356 10184
rect 39052 10060 39092 10100
rect 39340 10060 39380 10100
rect 43852 10060 43892 10100
rect 44428 10060 44468 10100
rect 46348 10060 46388 10100
rect 46732 10060 46772 10100
rect 49900 10060 49940 10100
rect 53068 10060 53108 10100
rect 53644 10060 53684 10100
rect 59212 10060 59252 10100
rect 64684 10060 64724 10100
rect 68812 10060 68852 10100
rect 70444 10060 70484 10100
rect 73420 10060 73460 10100
rect 77068 10060 77108 10100
rect 652 9976 692 10016
rect 42316 9976 42356 10016
rect 52300 9976 52340 10016
rect 58348 9976 58388 10016
rect 59692 9976 59732 10016
rect 59884 9976 59924 10016
rect 75820 9976 75860 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 1516 9640 1556 9680
rect 7180 9640 7220 9680
rect 40108 9640 40148 9680
rect 52684 9640 52724 9680
rect 53068 9640 53108 9680
rect 61996 9640 62036 9680
rect 64588 9640 64628 9680
rect 69292 9640 69332 9680
rect 69676 9640 69716 9680
rect 75532 9640 75572 9680
rect 77164 9640 77204 9680
rect 4492 9556 4532 9596
rect 4780 9556 4820 9596
rect 62188 9556 62228 9596
rect 64876 9556 64916 9596
rect 65356 9556 65396 9596
rect 66892 9556 66932 9596
rect 1996 9472 2036 9512
rect 2092 9472 2132 9512
rect 2188 9472 2228 9512
rect 2284 9472 2324 9512
rect 2860 9487 2900 9527
rect 3148 9472 3188 9512
rect 3244 9472 3284 9512
rect 3724 9472 3764 9512
rect 3916 9472 3956 9512
rect 4300 9472 4340 9512
rect 4396 9472 4436 9512
rect 4588 9472 4628 9512
rect 5164 9472 5204 9512
rect 6028 9472 6068 9512
rect 39148 9472 39188 9512
rect 39244 9472 39284 9512
rect 39436 9472 39476 9512
rect 39916 9472 39956 9512
rect 40012 9472 40052 9512
rect 40204 9472 40244 9512
rect 40588 9472 40628 9512
rect 40684 9472 40724 9512
rect 40780 9472 40820 9512
rect 40876 9472 40916 9512
rect 41644 9472 41684 9512
rect 41740 9472 41780 9512
rect 41932 9472 41972 9512
rect 42124 9472 42164 9512
rect 42220 9472 42260 9512
rect 42412 9472 42452 9512
rect 42604 9472 42644 9512
rect 42700 9472 42740 9512
rect 42796 9472 42836 9512
rect 42892 9472 42932 9512
rect 45868 9472 45908 9512
rect 46060 9472 46100 9512
rect 46540 9472 46580 9512
rect 46636 9472 46676 9512
rect 46924 9472 46964 9512
rect 50668 9472 50708 9512
rect 52972 9472 53012 9512
rect 53164 9472 53204 9512
rect 53270 9453 53310 9493
rect 53740 9472 53780 9512
rect 53932 9472 53972 9512
rect 54220 9472 54260 9512
rect 54412 9472 54452 9512
rect 57772 9472 57812 9512
rect 57964 9472 58004 9512
rect 58060 9472 58100 9512
rect 58348 9472 58388 9512
rect 58636 9472 58676 9512
rect 58732 9472 58772 9512
rect 59596 9472 59636 9512
rect 59980 9472 60020 9512
rect 60844 9472 60884 9512
rect 62572 9472 62612 9512
rect 63436 9472 63476 9512
rect 64780 9472 64820 9512
rect 64972 9472 65012 9512
rect 65068 9472 65108 9512
rect 65260 9472 65300 9512
rect 65452 9472 65492 9512
rect 67276 9472 67316 9512
rect 68140 9472 68180 9512
rect 69868 9472 69908 9512
rect 70060 9472 70100 9512
rect 70156 9472 70196 9512
rect 70732 9472 70772 9512
rect 70828 9472 70868 9512
rect 70924 9472 70964 9512
rect 71308 9472 71348 9512
rect 71500 9472 71540 9512
rect 71692 9472 71732 9512
rect 71884 9472 71924 9512
rect 75628 9472 75668 9512
rect 75724 9493 75764 9533
rect 75820 9493 75860 9533
rect 76012 9472 76052 9512
rect 76204 9485 76244 9525
rect 76300 9472 76340 9512
rect 77068 9472 77108 9512
rect 77260 9472 77300 9512
rect 77356 9472 77396 9512
rect 77548 9472 77588 9512
rect 77740 9472 77780 9512
rect 77932 9472 77972 9512
rect 78124 9472 78164 9512
rect 844 9388 884 9428
rect 1708 9388 1748 9428
rect 52108 9388 52148 9428
rect 57388 9388 57428 9428
rect 59404 9388 59444 9428
rect 3532 9346 3572 9386
rect 69474 9385 69514 9425
rect 70348 9388 70388 9428
rect 76492 9388 76532 9428
rect 1324 9304 1364 9344
rect 39436 9304 39476 9344
rect 41452 9304 41492 9344
rect 41932 9304 41972 9344
rect 44716 9304 44756 9344
rect 46252 9304 46292 9344
rect 47212 9304 47252 9344
rect 50380 9304 50420 9344
rect 54892 9304 54932 9344
rect 56428 9304 56468 9344
rect 69868 9304 69908 9344
rect 72172 9304 72212 9344
rect 73900 9304 73940 9344
rect 76012 9304 76052 9344
rect 77644 9304 77684 9344
rect 652 9220 692 9260
rect 3820 9220 3860 9260
rect 7180 9220 7220 9260
rect 42412 9220 42452 9260
rect 45964 9220 46004 9260
rect 52684 9220 52724 9260
rect 53836 9220 53876 9260
rect 54316 9220 54356 9260
rect 57580 9220 57620 9260
rect 57772 9220 57812 9260
rect 59020 9220 59060 9260
rect 59212 9220 59252 9260
rect 61996 9220 62036 9260
rect 64588 9220 64628 9260
rect 69292 9220 69332 9260
rect 69676 9220 69716 9260
rect 70540 9220 70580 9260
rect 71404 9220 71444 9260
rect 71788 9220 71828 9260
rect 76684 9220 76724 9260
rect 78028 9220 78068 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 43948 8884 43988 8924
rect 46636 8884 46676 8924
rect 51340 8884 51380 8924
rect 53932 8884 53972 8924
rect 56812 8884 56852 8924
rect 69772 8884 69812 8924
rect 71500 8884 71540 8924
rect 74092 8884 74132 8924
rect 79468 8884 79508 8924
rect 49324 8800 49364 8840
rect 844 8716 884 8756
rect 3532 8716 3572 8756
rect 50956 8758 50996 8798
rect 58924 8800 58964 8840
rect 60940 8800 60980 8840
rect 66508 8800 66548 8840
rect 68524 8800 68564 8840
rect 69196 8800 69236 8840
rect 70060 8800 70100 8840
rect 74284 8800 74324 8840
rect 76876 8800 76916 8840
rect 58252 8716 58292 8756
rect 58732 8716 58772 8756
rect 59692 8716 59732 8756
rect 64780 8716 64820 8756
rect 70252 8716 70292 8756
rect 1516 8632 1556 8672
rect 2380 8632 2420 8672
rect 4780 8632 4820 8672
rect 4972 8632 5012 8672
rect 41932 8632 41972 8672
rect 42796 8632 42836 8672
rect 44620 8632 44660 8672
rect 45484 8632 45524 8672
rect 48460 8632 48500 8672
rect 48652 8632 48692 8672
rect 48844 8632 48884 8672
rect 49036 8632 49076 8672
rect 49132 8632 49172 8672
rect 49708 8632 49748 8672
rect 49804 8632 49844 8672
rect 49900 8632 49940 8672
rect 51340 8632 51380 8672
rect 51532 8632 51572 8672
rect 51628 8632 51668 8672
rect 52204 8632 52244 8672
rect 52300 8632 52340 8672
rect 52396 8632 52436 8672
rect 52492 8632 52532 8672
rect 52684 8632 52724 8672
rect 52876 8632 52916 8672
rect 52972 8632 53012 8672
rect 53260 8649 53300 8689
rect 53548 8632 53588 8672
rect 54796 8632 54836 8672
rect 55660 8632 55700 8672
rect 57772 8632 57812 8672
rect 57868 8632 57908 8672
rect 57964 8632 58004 8672
rect 58060 8632 58100 8672
rect 59116 8632 59156 8672
rect 59308 8632 59348 8672
rect 59404 8632 59444 8672
rect 59596 8632 59636 8672
rect 59788 8632 59828 8672
rect 59980 8632 60020 8672
rect 60076 8632 60116 8672
rect 60172 8632 60212 8672
rect 63820 8632 63860 8672
rect 63916 8632 63956 8672
rect 64012 8632 64052 8672
rect 64108 8632 64148 8672
rect 64300 8632 64340 8672
rect 64492 8632 64532 8672
rect 64588 8632 64628 8672
rect 68716 8632 68756 8672
rect 68908 8632 68948 8672
rect 69004 8632 69044 8672
rect 69196 8632 69236 8672
rect 69388 8632 69428 8672
rect 69484 8632 69524 8672
rect 69676 8611 69716 8651
rect 69868 8632 69908 8672
rect 70828 8632 70868 8672
rect 71116 8632 71156 8672
rect 72076 8632 72116 8672
rect 72940 8632 72980 8672
rect 75628 8632 75668 8672
rect 75820 8632 75860 8672
rect 75916 8632 75956 8672
rect 76204 8632 76244 8672
rect 76492 8632 76532 8672
rect 77452 8632 77492 8672
rect 78316 8632 78356 8672
rect 1132 8548 1172 8588
rect 4876 8548 4916 8588
rect 41548 8548 41588 8588
rect 44236 8548 44276 8588
rect 48556 8548 48596 8588
rect 53644 8548 53684 8588
rect 54412 8548 54452 8588
rect 59212 8548 59252 8588
rect 64396 8548 64436 8588
rect 71212 8548 71252 8588
rect 71692 8548 71732 8588
rect 75724 8548 75764 8588
rect 76588 8548 76628 8588
rect 77068 8548 77108 8588
rect 652 8464 692 8504
rect 43948 8464 43988 8504
rect 46636 8464 46676 8504
rect 48940 8464 48980 8504
rect 52780 8464 52820 8504
rect 58444 8464 58484 8504
rect 64972 8464 65012 8504
rect 68812 8464 68852 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 2380 8128 2420 8168
rect 4684 8128 4724 8168
rect 7468 8128 7508 8168
rect 45004 8128 45044 8168
rect 52876 8128 52916 8168
rect 58348 8128 58388 8168
rect 62860 8128 62900 8168
rect 64108 8128 64148 8168
rect 65644 8128 65684 8168
rect 68428 8128 68468 8168
rect 71020 8128 71060 8168
rect 71500 8128 71540 8168
rect 75916 8128 75956 8168
rect 77068 8128 77108 8168
rect 5068 8044 5108 8084
rect 54124 8044 54164 8084
rect 55948 8044 55988 8084
rect 66028 8044 66068 8084
rect 68620 8044 68660 8084
rect 1804 7960 1844 8000
rect 1900 7960 1940 8000
rect 1996 7960 2036 8000
rect 2092 7960 2132 8000
rect 2284 7960 2324 8000
rect 2476 7960 2516 8000
rect 2572 7960 2612 8000
rect 2764 7960 2804 8000
rect 2956 7960 2996 8000
rect 3052 7960 3092 8000
rect 3436 7960 3476 8000
rect 3724 7960 3764 8000
rect 3820 7960 3860 8000
rect 4588 7960 4628 8000
rect 4780 7960 4820 8000
rect 4876 7960 4916 8000
rect 5452 7960 5492 8000
rect 6316 7960 6356 8000
rect 44140 7960 44180 8000
rect 44236 7960 44276 8000
rect 44428 7960 44468 8000
rect 44812 7960 44852 8000
rect 44908 7960 44948 8000
rect 45100 7960 45140 8000
rect 45388 7960 45428 8000
rect 45484 7960 45524 8000
rect 45580 7960 45620 8000
rect 45676 7960 45716 8000
rect 46732 7960 46772 8000
rect 46828 7960 46868 8000
rect 47020 7960 47060 8000
rect 47212 7960 47252 8000
rect 47308 7960 47348 8000
rect 47500 7960 47540 8000
rect 47980 7960 48020 8000
rect 48268 7960 48308 8000
rect 48364 7960 48404 8000
rect 48844 7959 48884 7999
rect 49228 7960 49268 8000
rect 50188 7960 50228 8000
rect 50476 7960 50516 8000
rect 50860 7960 50900 8000
rect 51724 7960 51764 8000
rect 53068 7960 53108 8000
rect 53164 7960 53204 8000
rect 53260 7981 53300 8021
rect 53356 7960 53396 8000
rect 54028 7960 54068 8000
rect 54220 7960 54260 8000
rect 54316 7960 54356 8000
rect 56332 7960 56372 8000
rect 57196 7960 57236 8000
rect 58540 7960 58580 8000
rect 58636 7960 58676 8000
rect 58828 7960 58868 8000
rect 60076 7960 60116 8000
rect 60268 7960 60308 8000
rect 60460 7960 60500 8000
rect 60844 7960 60884 8000
rect 61708 7960 61748 8000
rect 63628 7960 63668 8000
rect 63820 7960 63860 8000
rect 63916 7960 63956 8000
rect 64204 7960 64244 8000
rect 64300 7960 64340 8000
rect 64396 7960 64436 8000
rect 64684 7960 64724 8000
rect 64972 7960 65012 8000
rect 65068 7960 65108 8000
rect 65548 7960 65588 8000
rect 65740 7960 65780 8000
rect 65836 7960 65876 8000
rect 66412 7960 66452 8000
rect 67276 7960 67316 8000
rect 69004 7960 69044 8000
rect 69868 7960 69908 8000
rect 71404 7960 71444 8000
rect 71596 7960 71636 8000
rect 71692 7960 71732 8000
rect 73516 7960 73556 8000
rect 73900 7960 73940 8000
rect 74764 7960 74804 8000
rect 76108 7960 76148 8000
rect 76204 7960 76244 8000
rect 76300 7960 76340 8000
rect 76396 7960 76436 8000
rect 76588 7960 76628 8000
rect 76780 7960 76820 8000
rect 76972 7960 77012 8000
rect 77164 7960 77204 8000
rect 77260 7960 77300 8000
rect 844 7876 884 7916
rect 1228 7876 1268 7916
rect 1612 7792 1652 7832
rect 2764 7792 2804 7832
rect 44428 7792 44468 7832
rect 45868 7792 45908 7832
rect 47020 7792 47060 7832
rect 48652 7792 48692 7832
rect 63052 7792 63092 7832
rect 77740 7792 77780 7832
rect 652 7708 692 7748
rect 1036 7708 1076 7748
rect 4108 7708 4148 7748
rect 7468 7708 7508 7748
rect 47500 7708 47540 7748
rect 49900 7708 49940 7748
rect 58828 7708 58868 7748
rect 60172 7708 60212 7748
rect 63628 7708 63668 7748
rect 65356 7708 65396 7748
rect 68428 7708 68468 7748
rect 71020 7708 71060 7748
rect 76684 7708 76724 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 3916 7372 3956 7412
rect 5068 7372 5108 7412
rect 47788 7372 47828 7412
rect 51148 7372 51188 7412
rect 64588 7372 64628 7412
rect 65356 7372 65396 7412
rect 65932 7372 65972 7412
rect 75532 7372 75572 7412
rect 5548 7288 5588 7328
rect 51916 7288 51956 7328
rect 55084 7288 55124 7328
rect 69388 7288 69428 7328
rect 72460 7288 72500 7328
rect 77836 7288 77876 7328
rect 844 7204 884 7244
rect 54700 7204 54740 7244
rect 1900 7120 1940 7160
rect 2764 7120 2804 7160
rect 4204 7120 4244 7160
rect 4396 7120 4436 7160
rect 4972 7120 5012 7160
rect 5164 7120 5204 7160
rect 45388 7120 45428 7160
rect 45772 7120 45812 7160
rect 46636 7120 46676 7160
rect 48748 7120 48788 7160
rect 49132 7120 49172 7160
rect 49996 7120 50036 7160
rect 52780 7120 52820 7160
rect 52972 7120 53012 7160
rect 53068 7120 53108 7160
rect 1516 7036 1556 7076
rect 4300 7036 4340 7076
rect 52876 7036 52916 7076
rect 53260 7078 53300 7118
rect 53452 7120 53492 7160
rect 53548 7120 53588 7160
rect 54316 7120 54356 7160
rect 54508 7120 54548 7160
rect 57196 7120 57236 7160
rect 58060 7120 58100 7160
rect 59692 7120 59732 7160
rect 59980 7120 60020 7160
rect 60556 7120 60596 7160
rect 60652 7120 60692 7160
rect 60844 7120 60884 7160
rect 62188 7120 62228 7160
rect 62572 7120 62612 7160
rect 63436 7120 63476 7160
rect 64780 7120 64820 7160
rect 64972 7120 65012 7160
rect 65068 7120 65108 7160
rect 65260 7120 65300 7160
rect 65452 7120 65492 7160
rect 65836 7121 65876 7161
rect 66028 7120 66068 7160
rect 66220 7120 66260 7160
rect 66412 7120 66452 7160
rect 66604 7120 66644 7160
rect 66796 7120 66836 7160
rect 69580 7120 69620 7160
rect 69676 7120 69716 7160
rect 69772 7120 69812 7160
rect 69868 7120 69908 7160
rect 70060 7120 70100 7160
rect 70252 7120 70292 7160
rect 70348 7120 70388 7160
rect 71692 7120 71732 7160
rect 71884 7120 71924 7160
rect 71980 7120 72020 7160
rect 75532 7120 75572 7160
rect 75724 7120 75764 7160
rect 75820 7120 75860 7160
rect 76012 7131 76052 7171
rect 76204 7120 76244 7160
rect 76300 7120 76340 7160
rect 76972 7120 77012 7160
rect 77164 7120 77204 7160
rect 77452 7120 77492 7160
rect 77644 7120 77684 7160
rect 53356 7036 53396 7076
rect 54412 7036 54452 7076
rect 56812 7036 56852 7076
rect 60076 7036 60116 7076
rect 60748 7036 60788 7076
rect 64876 7036 64916 7076
rect 66316 7036 66356 7076
rect 66700 7036 66740 7076
rect 76108 7036 76148 7076
rect 77068 7036 77108 7076
rect 77548 7036 77588 7076
rect 652 6952 692 6992
rect 54892 6952 54932 6992
rect 59212 6952 59252 6992
rect 70156 6952 70196 6992
rect 71788 6952 71828 6992
rect 60364 6910 60404 6950
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 2188 6616 2228 6656
rect 7468 6616 7508 6656
rect 47212 6616 47252 6656
rect 53836 6616 53876 6656
rect 57004 6616 57044 6656
rect 69004 6616 69044 6656
rect 74380 6616 74420 6656
rect 79468 6616 79508 6656
rect 54220 6532 54260 6572
rect 54604 6532 54644 6572
rect 66028 6532 66068 6572
rect 71980 6532 72020 6572
rect 2092 6448 2132 6488
rect 2284 6448 2324 6488
rect 2380 6448 2420 6488
rect 2572 6448 2612 6488
rect 2764 6448 2804 6488
rect 2870 6429 2910 6469
rect 4108 6448 4148 6488
rect 4204 6448 4244 6488
rect 4492 6448 4532 6488
rect 5068 6448 5108 6488
rect 5452 6448 5492 6488
rect 6316 6448 6356 6488
rect 47308 6448 47348 6488
rect 47404 6448 47444 6488
rect 47500 6448 47540 6488
rect 47692 6448 47732 6488
rect 47884 6448 47924 6488
rect 47980 6448 48020 6488
rect 48364 6448 48404 6488
rect 48556 6448 48596 6488
rect 48844 6448 48884 6488
rect 49228 6448 49268 6488
rect 50092 6448 50132 6488
rect 51436 6448 51476 6488
rect 51820 6448 51860 6488
rect 52684 6448 52724 6488
rect 54124 6448 54164 6488
rect 54316 6448 54356 6488
rect 54412 6448 54452 6488
rect 54988 6448 55028 6488
rect 55852 6448 55892 6488
rect 58060 6448 58100 6488
rect 58252 6448 58292 6488
rect 58348 6448 58388 6488
rect 58540 6448 58580 6488
rect 58636 6448 58676 6488
rect 58732 6448 58772 6488
rect 58828 6448 58868 6488
rect 59212 6448 59252 6488
rect 59308 6448 59348 6488
rect 59500 6448 59540 6488
rect 60172 6448 60212 6488
rect 60364 6448 60404 6488
rect 61036 6448 61076 6488
rect 61228 6448 61268 6488
rect 61324 6448 61364 6488
rect 65644 6448 65684 6488
rect 65932 6448 65972 6488
rect 66604 6448 66644 6488
rect 66988 6448 67028 6488
rect 67852 6448 67892 6488
rect 69196 6448 69236 6488
rect 69580 6448 69620 6488
rect 70444 6448 70484 6488
rect 72364 6448 72404 6488
rect 73228 6448 73268 6488
rect 75628 6448 75668 6488
rect 75724 6448 75764 6488
rect 75820 6448 75860 6488
rect 75916 6448 75956 6488
rect 76204 6448 76244 6488
rect 76492 6448 76532 6488
rect 76588 6448 76628 6488
rect 77068 6448 77108 6488
rect 77452 6448 77492 6488
rect 78316 6448 78356 6488
rect 1708 6280 1748 6320
rect 2572 6280 2612 6320
rect 57292 6280 57332 6320
rect 58060 6280 58100 6320
rect 60268 6280 60308 6320
rect 61708 6280 61748 6320
rect 63436 6280 63476 6320
rect 66316 6280 66356 6320
rect 74764 6280 74804 6320
rect 76876 6280 76916 6320
rect 3820 6196 3860 6236
rect 47692 6196 47732 6236
rect 48460 6196 48500 6236
rect 51244 6196 51284 6236
rect 53836 6196 53876 6236
rect 57004 6196 57044 6236
rect 59500 6196 59540 6236
rect 61036 6196 61076 6236
rect 71596 6196 71636 6236
rect 74380 6196 74420 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 6316 5860 6356 5900
rect 48748 5860 48788 5900
rect 48940 5860 48980 5900
rect 54508 5860 54548 5900
rect 66316 5860 66356 5900
rect 69772 5860 69812 5900
rect 72652 5860 72692 5900
rect 73612 5860 73652 5900
rect 77164 5860 77204 5900
rect 46156 5776 46196 5816
rect 49420 5776 49460 5816
rect 56620 5776 56660 5816
rect 59692 5776 59732 5816
rect 61036 5776 61076 5816
rect 67180 5776 67220 5816
rect 71980 5776 72020 5816
rect 1036 5692 1076 5732
rect 3628 5692 3668 5732
rect 54796 5692 54836 5732
rect 1612 5608 1652 5648
rect 2476 5608 2516 5648
rect 5740 5608 5780 5648
rect 6028 5608 6068 5648
rect 6124 5608 6164 5648
rect 6316 5608 6356 5648
rect 47212 5608 47252 5648
rect 47404 5608 47444 5648
rect 47500 5608 47540 5648
rect 48076 5608 48116 5648
rect 48364 5608 48404 5648
rect 48940 5608 48980 5648
rect 49132 5608 49172 5648
rect 49228 5608 49268 5648
rect 52204 5608 52244 5648
rect 52300 5608 52340 5648
rect 52492 5608 52532 5648
rect 52780 5608 52820 5648
rect 52876 5608 52916 5648
rect 52972 5608 53012 5648
rect 53836 5608 53876 5648
rect 54124 5608 54164 5648
rect 54220 5608 54260 5648
rect 54700 5608 54740 5648
rect 54892 5608 54932 5648
rect 56236 5608 56276 5648
rect 56428 5608 56468 5648
rect 59212 5608 59252 5648
rect 59404 5608 59444 5648
rect 59500 5608 59540 5648
rect 60364 5608 60404 5648
rect 60652 5608 60692 5648
rect 61228 5608 61268 5648
rect 61612 5608 61652 5648
rect 62476 5608 62516 5648
rect 64588 5608 64628 5648
rect 64780 5608 64820 5648
rect 64876 5608 64916 5648
rect 65068 5608 65108 5648
rect 65164 5608 65204 5648
rect 65260 5608 65300 5648
rect 65356 5608 65396 5648
rect 1228 5524 1268 5564
rect 48460 5524 48500 5564
rect 52396 5524 52436 5564
rect 52684 5524 52724 5564
rect 56332 5524 56372 5564
rect 60748 5524 60788 5564
rect 66316 5566 66356 5606
rect 66508 5608 66548 5648
rect 66604 5608 66644 5648
rect 69292 5587 69332 5627
rect 69388 5608 69428 5648
rect 69484 5608 69524 5648
rect 69580 5608 69620 5648
rect 69772 5608 69812 5648
rect 69964 5608 70004 5648
rect 70060 5608 70100 5648
rect 71308 5608 71348 5648
rect 71596 5608 71636 5648
rect 71692 5608 71732 5648
rect 72172 5608 72212 5648
rect 72364 5608 72404 5648
rect 72556 5608 72596 5648
rect 72748 5608 72788 5648
rect 74764 5608 74804 5648
rect 75628 5608 75668 5648
rect 76204 5608 76244 5648
rect 76396 5608 76436 5648
rect 76492 5608 76532 5648
rect 77164 5608 77204 5648
rect 77356 5608 77396 5648
rect 77452 5608 77492 5648
rect 72268 5524 72308 5564
rect 76012 5524 76052 5564
rect 844 5440 884 5480
rect 47308 5440 47348 5480
rect 59308 5440 59348 5480
rect 63628 5440 63668 5480
rect 64684 5440 64724 5480
rect 76300 5440 76340 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 652 5104 692 5144
rect 2188 5104 2228 5144
rect 52204 5104 52244 5144
rect 55756 5104 55796 5144
rect 65356 5104 65396 5144
rect 65644 5104 65684 5144
rect 76108 5104 76148 5144
rect 3532 5020 3572 5060
rect 3916 5020 3956 5060
rect 4300 5020 4340 5060
rect 45676 5020 45716 5060
rect 48556 5020 48596 5060
rect 52588 5020 52628 5060
rect 56140 5020 56180 5060
rect 58828 5020 58868 5060
rect 61900 5020 61940 5060
rect 62956 5020 62996 5060
rect 1612 4936 1652 4976
rect 1708 4936 1748 4976
rect 1804 4936 1844 4976
rect 1900 4936 1940 4976
rect 2092 4936 2132 4976
rect 2284 4936 2324 4976
rect 2380 4936 2420 4976
rect 3436 4936 3476 4976
rect 3628 4936 3668 4976
rect 3820 4936 3860 4976
rect 4012 4936 4052 4976
rect 5164 4936 5204 4976
rect 46060 4936 46100 4976
rect 46924 4936 46964 4976
rect 48460 4936 48500 4976
rect 48652 4936 48692 4976
rect 48844 4936 48884 4976
rect 48940 4936 48980 4976
rect 49132 4936 49172 4976
rect 51532 4936 51572 4976
rect 51724 4936 51764 4976
rect 51820 4936 51860 4976
rect 52012 4936 52052 4976
rect 52108 4936 52148 4976
rect 52300 4936 52340 4976
rect 52492 4936 52532 4976
rect 52684 4936 52724 4976
rect 55660 4936 55700 4976
rect 55852 4936 55892 4976
rect 55948 4936 55988 4976
rect 56524 4936 56564 4976
rect 57388 4936 57428 4976
rect 59212 4936 59252 4976
rect 60076 4936 60116 4976
rect 61420 4936 61460 4976
rect 61612 4936 61652 4976
rect 61804 4936 61844 4976
rect 61996 4936 62036 4976
rect 63340 4936 63380 4976
rect 64204 4936 64244 4976
rect 65548 4936 65588 4976
rect 65740 4936 65780 4976
rect 65836 4936 65876 4976
rect 66124 4936 66164 4976
rect 66316 4936 66356 4976
rect 66508 4936 66548 4976
rect 66700 4936 66740 4976
rect 68812 4936 68852 4976
rect 69004 4936 69044 4976
rect 69100 4936 69140 4976
rect 71212 4936 71252 4976
rect 71404 4936 71444 4976
rect 71596 4936 71636 4976
rect 71788 4936 71828 4976
rect 71884 4936 71924 4976
rect 75916 4936 75956 4976
rect 76012 4936 76052 4976
rect 76204 4936 76244 4976
rect 76396 4936 76436 4976
rect 76588 4936 76628 4976
rect 76684 4936 76724 4976
rect 77164 4936 77204 4976
rect 77356 4936 77396 4976
rect 77452 4936 77492 4976
rect 844 4852 884 4892
rect 1420 4852 1460 4892
rect 5548 4768 5588 4808
rect 5932 4768 5972 4808
rect 50092 4768 50132 4808
rect 52876 4768 52916 4808
rect 61516 4768 61556 4808
rect 66892 4768 66932 4808
rect 69484 4768 69524 4808
rect 72364 4768 72404 4808
rect 74476 4768 74516 4808
rect 77836 4768 77876 4808
rect 1228 4684 1268 4724
rect 48076 4684 48116 4724
rect 49132 4684 49172 4724
rect 51532 4684 51572 4724
rect 58540 4684 58580 4724
rect 61228 4684 61268 4724
rect 66220 4684 66260 4724
rect 66604 4684 66644 4724
rect 68812 4684 68852 4724
rect 71308 4684 71348 4724
rect 71596 4684 71636 4724
rect 76396 4684 76436 4724
rect 77164 4684 77204 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 2380 4348 2420 4388
rect 52012 4348 52052 4388
rect 66220 4348 66260 4388
rect 652 4264 692 4304
rect 1804 4264 1844 4304
rect 4204 4264 4244 4304
rect 5068 4264 5108 4304
rect 7660 4264 7700 4304
rect 54700 4264 54740 4304
rect 55084 4264 55124 4304
rect 56812 4264 56852 4304
rect 57964 4264 58004 4304
rect 60172 4264 60212 4304
rect 68812 4264 68852 4304
rect 74284 4264 74324 4304
rect 76876 4264 76916 4304
rect 79468 4264 79508 4304
rect 844 4180 884 4220
rect 1228 4180 1268 4220
rect 4492 4180 4532 4220
rect 2380 4096 2420 4136
rect 2572 4096 2612 4136
rect 2668 4096 2708 4136
rect 2860 4054 2900 4094
rect 3052 4096 3092 4136
rect 3148 4096 3188 4136
rect 3532 4096 3572 4136
rect 3820 4096 3860 4136
rect 4396 4096 4436 4136
rect 4588 4096 4628 4136
rect 4780 4096 4820 4136
rect 4876 4096 4916 4136
rect 5068 4096 5108 4136
rect 5260 4096 5300 4136
rect 5644 4096 5684 4136
rect 6508 4096 6548 4136
rect 47404 4096 47444 4136
rect 47500 4096 47540 4136
rect 47596 4096 47636 4136
rect 47692 4096 47732 4136
rect 49996 4096 50036 4136
rect 50860 4096 50900 4136
rect 52300 4096 52340 4136
rect 52684 4096 52724 4136
rect 53548 4096 53588 4136
rect 55564 4096 55604 4136
rect 55660 4096 55700 4136
rect 55756 4096 55796 4136
rect 55852 4096 55892 4136
rect 56140 4096 56180 4136
rect 56428 4096 56468 4136
rect 57004 4096 57044 4136
rect 57196 4096 57236 4136
rect 57292 4096 57332 4136
rect 57964 4096 58004 4136
rect 58156 4096 58196 4136
rect 58252 4096 58292 4136
rect 58924 4096 58964 4136
rect 59020 4096 59060 4136
rect 59116 4096 59156 4136
rect 59212 4096 59252 4136
rect 63244 4096 63284 4136
rect 64108 4096 64148 4136
rect 65548 4096 65588 4136
rect 65836 4096 65876 4136
rect 66796 4096 66836 4136
rect 67660 4096 67700 4136
rect 69388 4096 69428 4136
rect 70252 4096 70292 4136
rect 71884 4096 71924 4136
rect 72268 4096 72308 4136
rect 73132 4096 73172 4136
rect 74476 4096 74516 4136
rect 74860 4096 74900 4136
rect 75724 4096 75764 4136
rect 77068 4096 77108 4136
rect 77452 4096 77492 4136
rect 78316 4096 78356 4136
rect 3916 4012 3956 4052
rect 49612 4012 49652 4052
rect 56524 4012 56564 4052
rect 62860 4012 62900 4052
rect 65932 4012 65972 4052
rect 66412 4012 66452 4052
rect 69004 4012 69044 4052
rect 1036 3928 1076 3968
rect 2956 3928 2996 3968
rect 52012 3928 52052 3968
rect 57100 3928 57140 3968
rect 65260 3928 65300 3968
rect 71404 3928 71444 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 3724 3592 3764 3632
rect 50188 3592 50228 3632
rect 62092 3592 62132 3632
rect 64012 3592 64052 3632
rect 66220 3592 66260 3632
rect 69292 3592 69332 3632
rect 76108 3592 76148 3632
rect 1324 3508 1364 3548
rect 4396 3508 4436 3548
rect 52012 3508 52052 3548
rect 56140 3508 56180 3548
rect 56716 3508 56756 3548
rect 71404 3508 71444 3548
rect 72172 3508 72212 3548
rect 76780 3508 76820 3548
rect 77356 3508 77396 3548
rect 77740 3508 77780 3548
rect 1708 3424 1748 3464
rect 2572 3424 2612 3464
rect 4300 3424 4340 3464
rect 4492 3424 4532 3464
rect 49996 3424 50036 3464
rect 50092 3424 50132 3464
rect 50284 3424 50324 3464
rect 50572 3424 50612 3464
rect 50668 3424 50708 3464
rect 50764 3424 50804 3464
rect 50860 3424 50900 3464
rect 51628 3424 51668 3464
rect 51916 3424 51956 3464
rect 52492 3424 52532 3464
rect 52684 3424 52724 3464
rect 54892 3424 54932 3464
rect 55756 3424 55796 3464
rect 56620 3424 56660 3464
rect 56812 3424 56852 3464
rect 59308 3424 59348 3464
rect 59500 3424 59540 3464
rect 59692 3424 59732 3464
rect 60076 3424 60116 3464
rect 60940 3424 60980 3464
rect 63820 3424 63860 3464
rect 63916 3424 63956 3464
rect 64108 3424 64148 3464
rect 64300 3424 64340 3464
rect 64396 3424 64436 3464
rect 64492 3424 64532 3464
rect 64588 3424 64628 3464
rect 66124 3424 66164 3464
rect 66316 3424 66356 3464
rect 66412 3424 66452 3464
rect 68620 3424 68660 3464
rect 68716 3424 68756 3464
rect 68908 3424 68948 3464
rect 69100 3424 69140 3464
rect 69196 3424 69236 3464
rect 69388 3424 69428 3464
rect 69676 3424 69716 3464
rect 69772 3424 69812 3464
rect 69868 3424 69908 3464
rect 69964 3424 70004 3464
rect 70636 3424 70676 3464
rect 70732 3424 70772 3464
rect 70924 3424 70964 3464
rect 71500 3424 71540 3464
rect 71788 3424 71828 3464
rect 72076 3424 72116 3464
rect 72268 3424 72308 3464
rect 72460 3424 72500 3464
rect 72844 3424 72884 3464
rect 73036 3424 73076 3464
rect 75820 3424 75860 3464
rect 75916 3424 75956 3464
rect 76012 3424 76052 3464
rect 76396 3424 76436 3464
rect 76684 3424 76724 3464
rect 77260 3424 77300 3464
rect 77452 3424 77492 3464
rect 77644 3424 77684 3464
rect 77836 3424 77876 3464
rect 1132 3340 1172 3380
rect 52300 3256 52340 3296
rect 52588 3256 52628 3296
rect 63340 3298 63380 3338
rect 68908 3256 68948 3296
rect 71116 3256 71156 3296
rect 77068 3256 77108 3296
rect 940 3172 980 3212
rect 53740 3172 53780 3212
rect 59404 3172 59444 3212
rect 70924 3172 70964 3212
rect 72940 3172 72980 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 652 2836 692 2876
rect 3052 2836 3092 2876
rect 58828 2836 58868 2876
rect 64012 2836 64052 2876
rect 72652 2836 72692 2876
rect 73324 2836 73364 2876
rect 76204 2836 76244 2876
rect 1516 2752 1556 2792
rect 53932 2752 53972 2792
rect 56908 2752 56948 2792
rect 60076 2752 60116 2792
rect 62188 2752 62228 2792
rect 66508 2752 66548 2792
rect 68716 2752 68756 2792
rect 70924 2752 70964 2792
rect 74668 2752 74708 2792
rect 76012 2752 76052 2792
rect 77452 2752 77492 2792
rect 78220 2752 78260 2792
rect 844 2668 884 2708
rect 1228 2668 1268 2708
rect 1708 2668 1748 2708
rect 60364 2668 60404 2708
rect 64780 2668 64820 2708
rect 2476 2584 2516 2624
rect 2572 2584 2612 2624
rect 2668 2584 2708 2624
rect 2764 2584 2804 2624
rect 3052 2584 3092 2624
rect 3244 2584 3284 2624
rect 3340 2584 3380 2624
rect 55756 2584 55796 2624
rect 55852 2584 55892 2624
rect 56044 2542 56084 2582
rect 56332 2584 56372 2624
rect 56524 2584 56564 2624
rect 56620 2584 56660 2624
rect 56812 2584 56852 2624
rect 57004 2584 57044 2624
rect 57196 2584 57236 2624
rect 57292 2584 57332 2624
rect 57484 2584 57524 2624
rect 58828 2584 58868 2624
rect 59020 2584 59060 2624
rect 59116 2584 59156 2624
rect 59404 2584 59444 2624
rect 59692 2584 59732 2624
rect 60268 2584 60308 2624
rect 60460 2584 60500 2624
rect 63724 2584 63764 2624
rect 63820 2584 63860 2624
rect 64012 2584 64052 2624
rect 64204 2584 64244 2624
rect 64396 2584 64436 2624
rect 64492 2584 64532 2624
rect 64684 2584 64724 2624
rect 64876 2584 64916 2624
rect 68236 2584 68276 2624
rect 68332 2584 68372 2624
rect 68428 2584 68468 2624
rect 68620 2584 68660 2624
rect 68812 2584 68852 2624
rect 69004 2584 69044 2624
rect 69196 2584 69236 2624
rect 71116 2584 71156 2624
rect 71212 2584 71252 2624
rect 71404 2584 71444 2624
rect 71596 2584 71636 2624
rect 71692 2621 71732 2661
rect 71788 2626 71828 2666
rect 71884 2584 71924 2624
rect 72172 2584 72212 2624
rect 73612 2584 73652 2624
rect 73708 2584 73748 2624
rect 73996 2584 74036 2624
rect 74284 2584 74324 2624
rect 74476 2584 74516 2624
rect 76204 2584 76244 2624
rect 76396 2584 76436 2624
rect 76492 2584 76532 2624
rect 76780 2584 76820 2624
rect 77068 2584 77108 2624
rect 77644 2584 77684 2624
rect 77836 2584 77876 2624
rect 59788 2500 59828 2540
rect 69100 2500 69140 2540
rect 74380 2500 74420 2540
rect 77164 2500 77204 2540
rect 77740 2500 77780 2540
rect 1036 2416 1076 2456
rect 55948 2416 55988 2456
rect 56428 2416 56468 2456
rect 57388 2416 57428 2456
rect 64300 2416 64340 2456
rect 68140 2416 68180 2456
rect 71308 2416 71348 2456
rect 72652 2416 72692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 55852 2080 55892 2120
rect 61612 2080 61652 2120
rect 66892 2080 66932 2120
rect 71212 2080 71252 2120
rect 73804 2080 73844 2120
rect 56620 1996 56660 2036
rect 64492 1996 64532 2036
rect 71404 1996 71444 2036
rect 53452 1912 53492 1952
rect 53836 1912 53876 1952
rect 54700 1912 54740 1952
rect 56044 1912 56084 1952
rect 56236 1912 56276 1952
rect 56332 1912 56372 1952
rect 57004 1912 57044 1952
rect 57868 1912 57908 1952
rect 59212 1912 59252 1952
rect 59596 1912 59636 1952
rect 60460 1912 60500 1952
rect 61804 1912 61844 1952
rect 62188 1912 62228 1952
rect 63052 1912 63092 1952
rect 64876 1912 64916 1952
rect 65740 1912 65780 1952
rect 67372 1912 67412 1952
rect 67564 1912 67604 1952
rect 67660 1912 67700 1952
rect 67948 1912 67988 1952
rect 68236 1912 68276 1952
rect 68332 1912 68372 1952
rect 68812 1912 68852 1952
rect 69196 1912 69236 1952
rect 70060 1912 70100 1952
rect 71788 1912 71828 1952
rect 72652 1912 72692 1952
rect 73996 1912 74036 1952
rect 74188 1912 74228 1952
rect 74284 1912 74324 1952
rect 74572 1912 74612 1952
rect 74668 1912 74708 1952
rect 74860 1912 74900 1952
rect 75148 1912 75188 1952
rect 75244 1912 75284 1952
rect 75436 1912 75476 1952
rect 75628 1912 75668 1952
rect 76012 1912 76052 1952
rect 76876 1912 76916 1952
rect 78220 1912 78260 1952
rect 78412 1912 78452 1952
rect 78508 1912 78548 1952
rect 78700 1912 78740 1952
rect 78892 1912 78932 1952
rect 56044 1744 56084 1784
rect 68620 1744 68660 1784
rect 74860 1744 74900 1784
rect 75436 1744 75476 1784
rect 78796 1744 78836 1784
rect 59020 1660 59060 1700
rect 61612 1660 61652 1700
rect 64204 1660 64244 1700
rect 67372 1660 67412 1700
rect 73996 1660 74036 1700
rect 78028 1660 78068 1700
rect 78220 1660 78260 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 56812 1324 56852 1364
rect 58924 1324 58964 1364
rect 62476 1324 62516 1364
rect 68428 1324 68468 1364
rect 68908 1324 68948 1364
rect 70156 1324 70196 1364
rect 71884 1324 71924 1364
rect 75628 1324 75668 1364
rect 77068 1324 77108 1364
rect 57100 1240 57140 1280
rect 57388 1240 57428 1280
rect 60844 1240 60884 1280
rect 61996 1240 62036 1280
rect 64492 1240 64532 1280
rect 64780 1240 64820 1280
rect 65068 1240 65108 1280
rect 69388 1240 69428 1280
rect 55468 1072 55508 1112
rect 55564 1072 55604 1112
rect 55660 1072 55700 1112
rect 55756 1072 55796 1112
rect 56140 1072 56180 1112
rect 56428 1072 56468 1112
rect 56524 1072 56564 1112
rect 57004 1072 57044 1112
rect 57196 1072 57236 1112
rect 58636 1072 58676 1112
rect 58732 1072 58772 1112
rect 58924 1072 58964 1112
rect 59116 1072 59156 1112
rect 60076 1072 60116 1112
rect 60460 1072 60500 1112
rect 60556 1072 60596 1112
rect 60652 1072 60692 1112
rect 61708 1072 61748 1112
rect 61804 1072 61844 1112
rect 61996 1072 62036 1112
rect 62188 1072 62228 1112
rect 62284 1072 62324 1112
rect 62476 1072 62516 1112
rect 62668 1072 62708 1112
rect 62764 1072 62804 1112
rect 62860 1072 62900 1112
rect 62956 1072 62996 1112
rect 63820 1072 63860 1112
rect 64108 1072 64148 1112
rect 64684 1072 64724 1112
rect 64876 1072 64916 1112
rect 66028 1072 66068 1112
rect 66412 1072 66452 1112
rect 67276 1072 67316 1112
rect 68620 1072 68660 1112
rect 68716 1072 68756 1112
rect 68908 1072 68948 1112
rect 70732 1072 70772 1112
rect 71212 1072 71252 1112
rect 72556 1072 72596 1112
rect 73228 1072 73268 1112
rect 73612 1072 73652 1112
rect 74476 1072 74516 1112
rect 76012 1072 76052 1112
rect 76108 1072 76148 1112
rect 76204 1072 76244 1112
rect 78220 1072 78260 1112
rect 79084 1072 79124 1112
rect 79468 1072 79508 1112
rect 64204 988 64244 1028
rect 60364 904 60404 944
rect 75916 904 75956 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 63820 38368 64148 38408
rect 58060 38240 58100 38249
rect 58252 38240 58292 38249
rect 58100 38200 58196 38240
rect 58060 38191 58100 38200
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 57292 38156 57332 38167
rect 57292 38081 57332 38116
rect 57676 38156 57716 38165
rect 56428 38072 56468 38081
rect 844 37988 884 37997
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 844 37460 884 37948
rect 55947 37988 55989 37997
rect 55947 37948 55948 37988
rect 55988 37948 55989 37988
rect 55947 37939 55989 37948
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 54892 37568 54932 37577
rect 844 37420 980 37460
rect 652 26060 692 26069
rect 652 25817 692 26020
rect 843 25976 885 25985
rect 843 25936 844 25976
rect 884 25936 885 25976
rect 843 25927 885 25936
rect 844 25842 884 25927
rect 651 25808 693 25817
rect 651 25768 652 25808
rect 692 25768 693 25808
rect 651 25759 693 25768
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 844 25002 884 25087
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 844 24380 884 24389
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 844 23885 884 24340
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 843 23876 885 23885
rect 843 23836 844 23876
rect 884 23836 885 23876
rect 843 23827 885 23836
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 844 23490 884 23575
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 23036 692 23045
rect 556 22996 652 23036
rect 556 22457 596 22996
rect 652 22987 692 22996
rect 844 22868 884 22877
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 844 21617 884 22828
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 843 21608 885 21617
rect 843 21568 844 21608
rect 884 21568 885 21608
rect 843 21559 885 21568
rect 940 21449 980 37420
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 54411 36812 54453 36821
rect 54411 36772 54412 36812
rect 54452 36772 54453 36812
rect 54411 36763 54453 36772
rect 38667 36728 38709 36737
rect 38667 36688 38668 36728
rect 38708 36688 38709 36728
rect 38667 36679 38709 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 3819 30596 3861 30605
rect 3819 30556 3820 30596
rect 3860 30556 3861 30596
rect 3819 30547 3861 30556
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3820 27824 3860 30547
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 38476 29168 38516 29177
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 38476 28589 38516 29128
rect 38475 28580 38517 28589
rect 38475 28540 38476 28580
rect 38516 28540 38517 28580
rect 38475 28531 38517 28540
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 3820 27775 3860 27784
rect 37803 27740 37845 27749
rect 37803 27700 37804 27740
rect 37844 27700 37845 27740
rect 37803 27691 37845 27700
rect 3724 27656 3764 27665
rect 3628 27616 3724 27656
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 2763 25136 2805 25145
rect 2763 25096 2764 25136
rect 2804 25096 2805 25136
rect 2763 25087 2805 25096
rect 1803 24044 1845 24053
rect 1803 24004 1804 24044
rect 1844 24004 1845 24044
rect 1803 23995 1845 24004
rect 2187 24044 2229 24053
rect 2187 24004 2188 24044
rect 2228 24004 2229 24044
rect 2187 23995 2229 24004
rect 1804 23876 1844 23995
rect 2188 23910 2228 23995
rect 1804 23827 1844 23836
rect 1995 23876 2037 23885
rect 1995 23836 1996 23876
rect 2036 23836 2037 23876
rect 1995 23827 2037 23836
rect 1996 23742 2036 23827
rect 1419 23624 1461 23633
rect 1419 23584 1420 23624
rect 1460 23584 1461 23624
rect 1419 23575 1461 23584
rect 1612 23624 1652 23633
rect 1420 23129 1460 23575
rect 1515 23204 1557 23213
rect 1612 23204 1652 23584
rect 1515 23164 1516 23204
rect 1556 23164 1652 23204
rect 1515 23155 1557 23164
rect 1419 23120 1461 23129
rect 1419 23080 1420 23120
rect 1460 23080 1461 23120
rect 1419 23071 1461 23080
rect 1516 23120 1556 23155
rect 1420 22952 1460 23071
rect 1516 23069 1556 23080
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 1941 23120
rect 1899 23071 1941 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 1900 22986 1940 23071
rect 2092 22986 2132 23071
rect 1516 22952 1556 22961
rect 1420 22912 1516 22952
rect 1516 22903 1556 22912
rect 1708 22868 1748 22877
rect 1900 22868 1940 22877
rect 1748 22828 1844 22868
rect 1708 22819 1748 22828
rect 939 21440 981 21449
rect 939 21400 940 21440
rect 980 21400 981 21440
rect 939 21391 981 21400
rect 1707 21356 1749 21365
rect 1707 21316 1708 21356
rect 1748 21316 1749 21356
rect 1707 21307 1749 21316
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 1708 20012 1748 21307
rect 1804 20096 1844 22828
rect 1900 22373 1940 22828
rect 1899 22364 1941 22373
rect 1899 22324 1900 22364
rect 1940 22324 1941 22364
rect 1899 22315 1941 22324
rect 2667 21356 2709 21365
rect 2667 21316 2668 21356
rect 2708 21316 2709 21356
rect 2667 21307 2709 21316
rect 2668 21222 2708 21307
rect 1804 20056 2036 20096
rect 1708 19972 1844 20012
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 1707 17828 1749 17837
rect 1707 17788 1708 17828
rect 1748 17788 1749 17828
rect 1707 17779 1749 17788
rect 1708 17694 1748 17779
rect 1516 17576 1556 17585
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 1516 17300 1556 17536
rect 1516 17260 1652 17300
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 1516 16400 1556 16409
rect 652 15737 692 16360
rect 1420 16360 1516 16400
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 844 15485 884 15570
rect 1036 15560 1076 15569
rect 843 15476 885 15485
rect 843 15436 844 15476
rect 884 15436 885 15476
rect 843 15427 885 15436
rect 652 15308 692 15317
rect 692 15268 884 15308
rect 652 15259 692 15268
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 652 14754 692 14839
rect 844 14804 884 15268
rect 1036 14981 1076 15520
rect 1420 15560 1460 16360
rect 1516 16351 1556 16360
rect 1420 15511 1460 15520
rect 1035 14972 1077 14981
rect 1035 14932 1036 14972
rect 1076 14932 1077 14972
rect 1035 14923 1077 14932
rect 1612 14888 1652 17260
rect 1707 17240 1749 17249
rect 1707 17200 1708 17240
rect 1748 17200 1749 17240
rect 1707 17191 1749 17200
rect 1420 14848 1652 14888
rect 844 14755 884 14764
rect 1228 14804 1268 14813
rect 1036 14552 1076 14561
rect 1036 14057 1076 14512
rect 1132 14216 1172 14225
rect 1228 14216 1268 14764
rect 1172 14176 1268 14216
rect 1132 14167 1172 14176
rect 1035 14048 1077 14057
rect 1035 14008 1036 14048
rect 1076 14008 1077 14048
rect 1035 13999 1077 14008
rect 1323 13964 1365 13973
rect 1323 13924 1324 13964
rect 1364 13924 1365 13964
rect 1323 13915 1365 13924
rect 1324 13830 1364 13915
rect 747 13796 789 13805
rect 747 13756 748 13796
rect 788 13756 789 13796
rect 747 13747 789 13756
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 652 12234 692 12319
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 748 8756 788 13747
rect 1420 13544 1460 14848
rect 1515 14720 1557 14729
rect 1515 14680 1516 14720
rect 1556 14680 1557 14720
rect 1515 14671 1557 14680
rect 1612 14720 1652 14729
rect 1708 14720 1748 17191
rect 1804 14897 1844 19972
rect 1996 16316 2036 20056
rect 2475 17240 2517 17249
rect 2475 17200 2476 17240
rect 2516 17200 2517 17240
rect 2475 17191 2517 17200
rect 2476 17106 2516 17191
rect 2667 16988 2709 16997
rect 2667 16948 2668 16988
rect 2708 16948 2709 16988
rect 2667 16939 2709 16948
rect 2668 16854 2708 16939
rect 2379 16400 2421 16409
rect 2379 16360 2380 16400
rect 2420 16360 2421 16400
rect 2379 16351 2421 16360
rect 1996 16267 2036 16276
rect 2188 16064 2228 16075
rect 2188 15989 2228 16024
rect 2187 15980 2229 15989
rect 2187 15940 2188 15980
rect 2228 15940 2229 15980
rect 2187 15931 2229 15940
rect 2187 15728 2229 15737
rect 2187 15688 2188 15728
rect 2228 15688 2229 15728
rect 2187 15679 2229 15688
rect 1995 14972 2037 14981
rect 1995 14932 1996 14972
rect 2036 14932 2037 14972
rect 1995 14923 2037 14932
rect 1803 14888 1845 14897
rect 1803 14848 1804 14888
rect 1844 14848 1845 14888
rect 1803 14839 1845 14848
rect 1996 14838 2036 14923
rect 1516 13964 1556 14671
rect 1612 14309 1652 14680
rect 1707 14680 1708 14720
rect 1707 14671 1748 14680
rect 1804 14720 1844 14729
rect 1996 14720 2036 14729
rect 1844 14680 1996 14720
rect 1804 14671 1844 14680
rect 1996 14671 2036 14680
rect 2188 14720 2228 15679
rect 2284 15560 2324 15569
rect 2284 14888 2324 15520
rect 2380 14972 2420 16351
rect 2572 16316 2612 16325
rect 2572 16157 2612 16276
rect 2764 16316 2804 25087
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3628 23129 3668 27616
rect 3724 27607 3764 27616
rect 37804 27606 37844 27691
rect 38188 27656 38228 27665
rect 3820 27404 3860 27413
rect 3724 27364 3820 27380
rect 3724 27340 3860 27364
rect 3627 23120 3669 23129
rect 3627 23080 3628 23120
rect 3668 23080 3669 23120
rect 3627 23071 3669 23080
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3243 22364 3285 22373
rect 3243 22324 3244 22364
rect 3284 22324 3285 22364
rect 3243 22315 3285 22324
rect 3244 22230 3284 22315
rect 3436 22112 3476 22121
rect 3476 22072 3668 22112
rect 3436 22063 3476 22072
rect 3244 21785 3284 21870
rect 3243 21776 3285 21785
rect 3243 21736 3244 21776
rect 3284 21736 3285 21776
rect 3243 21727 3285 21736
rect 3051 21608 3093 21617
rect 3051 21568 3052 21608
rect 3092 21568 3093 21608
rect 3051 21559 3093 21568
rect 3148 21608 3188 21617
rect 3340 21608 3380 21617
rect 2860 21513 2900 21522
rect 3052 21474 3092 21559
rect 2860 21113 2900 21473
rect 3148 21449 3188 21568
rect 3244 21568 3340 21608
rect 3147 21440 3189 21449
rect 3147 21400 3148 21440
rect 3188 21400 3189 21440
rect 3147 21391 3189 21400
rect 3244 21365 3284 21568
rect 3340 21559 3380 21568
rect 3243 21356 3285 21365
rect 3243 21316 3244 21356
rect 3284 21316 3285 21356
rect 3243 21307 3285 21316
rect 3531 21356 3573 21365
rect 3531 21316 3532 21356
rect 3572 21316 3573 21356
rect 3531 21307 3573 21316
rect 3532 21222 3572 21307
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3628 21113 3668 22072
rect 3724 21524 3764 27340
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 35116 26984 35156 26993
rect 38188 26984 38228 27616
rect 38284 26984 38324 26993
rect 35156 26944 35636 26984
rect 38188 26944 38284 26984
rect 35020 26816 35060 26825
rect 34828 26776 35020 26816
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 33483 26228 33525 26237
rect 33483 26188 33484 26228
rect 33524 26188 33525 26228
rect 33483 26179 33525 26188
rect 34251 26228 34293 26237
rect 34251 26188 34252 26228
rect 34292 26188 34293 26228
rect 34251 26179 34293 26188
rect 32715 26144 32757 26153
rect 32715 26104 32716 26144
rect 32756 26104 32757 26144
rect 32715 26095 32757 26104
rect 33148 26144 33188 26153
rect 31947 25976 31989 25985
rect 31947 25936 31948 25976
rect 31988 25936 31989 25976
rect 31947 25927 31989 25936
rect 31948 25842 31988 25927
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 30316 25472 30356 25481
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 29835 24716 29877 24725
rect 29835 24676 29836 24716
rect 29876 24676 29877 24716
rect 29835 24667 29877 24676
rect 29836 24582 29876 24667
rect 30220 24632 30260 24641
rect 30316 24632 30356 25432
rect 32716 25472 32756 26095
rect 33148 25901 33188 26104
rect 33484 25985 33524 26179
rect 33963 26144 34005 26153
rect 33963 26104 33964 26144
rect 34004 26104 34005 26144
rect 33963 26095 34005 26104
rect 33964 26010 34004 26095
rect 33483 25976 33525 25985
rect 33483 25936 33484 25976
rect 33524 25936 33525 25976
rect 33483 25927 33525 25936
rect 33147 25892 33189 25901
rect 33147 25852 33148 25892
rect 33188 25852 33189 25892
rect 33147 25843 33189 25852
rect 32716 25423 32756 25432
rect 31948 25304 31988 25313
rect 30260 24592 30356 24632
rect 31084 24632 31124 24641
rect 30220 24583 30260 24592
rect 31084 24557 31124 24592
rect 31083 24548 31125 24557
rect 31083 24508 31084 24548
rect 31124 24508 31125 24548
rect 31083 24499 31125 24508
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 28684 23960 28724 23969
rect 28724 23920 28820 23960
rect 28684 23911 28724 23920
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 28203 23204 28245 23213
rect 28203 23164 28204 23204
rect 28244 23164 28245 23204
rect 28203 23155 28245 23164
rect 3819 23120 3861 23129
rect 3819 23080 3820 23120
rect 3860 23080 3861 23120
rect 3819 23071 3861 23080
rect 3724 21475 3764 21484
rect 2859 21104 2901 21113
rect 2859 21064 2860 21104
rect 2900 21064 2901 21104
rect 2859 21055 2901 21064
rect 3627 21104 3669 21113
rect 3627 21064 3628 21104
rect 3668 21064 3669 21104
rect 3627 21055 3669 21064
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3820 18089 3860 23071
rect 28204 23070 28244 23155
rect 28588 23120 28628 23129
rect 28780 23120 28820 23920
rect 29547 23876 29589 23885
rect 29547 23836 29548 23876
rect 29588 23836 29589 23876
rect 29547 23827 29589 23836
rect 29452 23120 29492 23129
rect 28628 23080 28820 23120
rect 29260 23080 29452 23120
rect 28588 23071 28628 23080
rect 22059 23036 22101 23045
rect 22059 22996 22060 23036
rect 22100 22996 22101 23036
rect 22059 22987 22101 22996
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 5740 21524 5780 21533
rect 5547 21440 5589 21449
rect 5547 21400 5548 21440
rect 5588 21400 5589 21440
rect 5547 21391 5589 21400
rect 4779 21356 4821 21365
rect 4779 21316 4780 21356
rect 4820 21316 4821 21356
rect 4779 21307 4821 21316
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4780 18425 4820 21307
rect 5452 20768 5492 20777
rect 5548 20768 5588 21391
rect 5740 21365 5780 21484
rect 5931 21524 5973 21533
rect 5931 21484 5932 21524
rect 5972 21484 5973 21524
rect 5931 21475 5973 21484
rect 5932 21390 5972 21475
rect 5739 21356 5781 21365
rect 5739 21316 5740 21356
rect 5780 21316 5781 21356
rect 5739 21307 5781 21316
rect 6123 21356 6165 21365
rect 6123 21316 6124 21356
rect 6164 21316 6165 21356
rect 6123 21307 6165 21316
rect 6124 20777 6164 21307
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 5492 20728 5588 20768
rect 6123 20768 6165 20777
rect 6123 20728 6124 20768
rect 6164 20728 6165 20768
rect 4779 18416 4821 18425
rect 4779 18376 4780 18416
rect 4820 18376 4821 18416
rect 4779 18367 4821 18376
rect 3915 18164 3957 18173
rect 3915 18124 3916 18164
rect 3956 18124 3957 18164
rect 3915 18115 3957 18124
rect 3819 18080 3861 18089
rect 3819 18040 3820 18080
rect 3860 18040 3861 18080
rect 3819 18031 3861 18040
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 2764 16267 2804 16276
rect 3340 16232 3380 16241
rect 2571 16148 2613 16157
rect 2571 16108 2572 16148
rect 2612 16108 2613 16148
rect 2571 16099 2613 16108
rect 2955 16148 2997 16157
rect 2955 16108 2956 16148
rect 2996 16108 2997 16148
rect 2955 16099 2997 16108
rect 2956 16064 2996 16099
rect 2956 16013 2996 16024
rect 2667 15980 2709 15989
rect 2667 15940 2668 15980
rect 2708 15940 2709 15980
rect 2667 15931 2709 15940
rect 2380 14932 2612 14972
rect 2284 14848 2516 14888
rect 2188 14671 2228 14680
rect 2284 14720 2324 14729
rect 1707 14552 1747 14671
rect 1707 14512 1748 14552
rect 1611 14300 1653 14309
rect 1611 14260 1612 14300
rect 1652 14260 1653 14300
rect 1611 14251 1653 14260
rect 1708 14132 1748 14512
rect 2187 14300 2229 14309
rect 2187 14260 2188 14300
rect 2228 14260 2229 14300
rect 2187 14251 2229 14260
rect 1708 14092 1844 14132
rect 1708 13964 1748 13973
rect 1516 13924 1708 13964
rect 1708 13915 1748 13924
rect 1515 13796 1557 13805
rect 1515 13756 1516 13796
rect 1556 13756 1557 13796
rect 1515 13747 1557 13756
rect 1516 13662 1556 13747
rect 1420 13504 1556 13544
rect 1228 13376 1268 13385
rect 844 13336 1228 13376
rect 844 13292 884 13336
rect 1228 13327 1268 13336
rect 844 13243 884 13252
rect 1420 13292 1460 13301
rect 1420 13049 1460 13252
rect 1419 13040 1461 13049
rect 1419 13000 1420 13040
rect 1460 13000 1461 13040
rect 1419 12991 1461 13000
rect 1516 12536 1556 13504
rect 1420 12496 1556 12536
rect 1612 13208 1652 13217
rect 844 12452 884 12461
rect 844 12368 884 12412
rect 1323 12452 1365 12461
rect 1323 12412 1324 12452
rect 1364 12412 1365 12452
rect 1323 12403 1365 12412
rect 1132 12368 1172 12377
rect 844 12328 1132 12368
rect 1132 12319 1172 12328
rect 1324 12318 1364 12403
rect 1323 12200 1365 12209
rect 1323 12160 1324 12200
rect 1364 12160 1365 12200
rect 1323 12151 1365 12160
rect 1228 11864 1268 11873
rect 844 11824 1228 11864
rect 844 11780 884 11824
rect 1228 11815 1268 11824
rect 844 11731 884 11740
rect 1324 11108 1364 12151
rect 1420 12116 1460 12496
rect 1516 12293 1556 12378
rect 1612 12377 1652 13168
rect 1707 13208 1749 13217
rect 1707 13168 1708 13208
rect 1748 13168 1749 13208
rect 1707 13159 1749 13168
rect 1708 13074 1748 13159
rect 1804 12536 1844 14092
rect 1900 13376 1940 13385
rect 1940 13336 2132 13376
rect 1900 13327 1940 13336
rect 1900 13208 1940 13217
rect 1900 12704 1940 13168
rect 2092 13208 2132 13336
rect 2092 13159 2132 13168
rect 2188 13040 2228 14251
rect 2284 14225 2324 14680
rect 2379 14300 2421 14309
rect 2379 14260 2380 14300
rect 2420 14260 2421 14300
rect 2379 14251 2421 14260
rect 2283 14216 2325 14225
rect 2283 14176 2284 14216
rect 2324 14176 2325 14216
rect 2283 14167 2325 14176
rect 2380 14216 2420 14251
rect 2380 14165 2420 14176
rect 2379 13544 2421 13553
rect 2379 13504 2380 13544
rect 2420 13504 2421 13544
rect 2379 13495 2421 13504
rect 1900 12655 1940 12664
rect 2092 13000 2228 13040
rect 2092 12629 2132 13000
rect 2091 12620 2133 12629
rect 2091 12580 2092 12620
rect 2132 12580 2133 12620
rect 2091 12571 2133 12580
rect 1996 12557 2036 12566
rect 1804 12517 1996 12536
rect 1804 12496 2036 12517
rect 2092 12557 2132 12571
rect 2092 12508 2132 12517
rect 2380 12536 2420 13495
rect 2476 13385 2516 14848
rect 2572 14720 2612 14932
rect 2572 14671 2612 14680
rect 2572 13964 2612 13973
rect 2668 13964 2708 15931
rect 3340 15560 3380 16192
rect 3532 16232 3572 16241
rect 3572 16192 3668 16232
rect 3532 16183 3572 16192
rect 3436 16148 3476 16157
rect 3436 15737 3476 16108
rect 3628 16073 3668 16192
rect 3627 16064 3669 16073
rect 3627 16024 3628 16064
rect 3668 16024 3669 16064
rect 3627 16015 3669 16024
rect 3435 15728 3477 15737
rect 3435 15688 3436 15728
rect 3476 15688 3477 15728
rect 3435 15679 3477 15688
rect 3628 15728 3668 16015
rect 3628 15679 3668 15688
rect 3340 15520 3572 15560
rect 3436 15317 3476 15402
rect 2955 15308 2997 15317
rect 2955 15268 2956 15308
rect 2996 15268 2997 15308
rect 2955 15259 2997 15268
rect 3435 15308 3477 15317
rect 3435 15268 3436 15308
rect 3476 15268 3477 15308
rect 3435 15259 3477 15268
rect 2859 15140 2901 15149
rect 2859 15100 2860 15140
rect 2900 15100 2901 15140
rect 2859 15091 2901 15100
rect 2763 14888 2805 14897
rect 2763 14848 2764 14888
rect 2804 14848 2805 14888
rect 2763 14839 2805 14848
rect 2612 13924 2708 13964
rect 2764 14048 2804 14839
rect 2860 14762 2900 15091
rect 2956 14729 2996 15259
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3244 14972 3284 14981
rect 3532 14972 3572 15520
rect 3820 15476 3860 18031
rect 3820 15427 3860 15436
rect 3628 15308 3668 15317
rect 3668 15268 3860 15308
rect 3628 15259 3668 15268
rect 3284 14932 3572 14972
rect 3244 14923 3284 14932
rect 2860 14713 2900 14722
rect 2955 14720 2997 14729
rect 2955 14680 2956 14720
rect 2996 14680 2997 14720
rect 2955 14671 2997 14680
rect 2956 14586 2996 14671
rect 2955 14468 2997 14477
rect 2955 14428 2956 14468
rect 2996 14428 2997 14468
rect 2955 14419 2997 14428
rect 2859 14216 2901 14225
rect 2859 14176 2860 14216
rect 2900 14176 2901 14216
rect 2859 14167 2901 14176
rect 2860 14082 2900 14167
rect 2572 13915 2612 13924
rect 2764 13553 2804 14008
rect 2956 14048 2996 14419
rect 2763 13544 2805 13553
rect 2763 13504 2764 13544
rect 2804 13504 2900 13544
rect 2763 13495 2805 13504
rect 2475 13376 2517 13385
rect 2475 13336 2476 13376
rect 2516 13336 2517 13376
rect 2475 13327 2517 13336
rect 2763 13376 2805 13385
rect 2763 13336 2764 13376
rect 2804 13336 2805 13376
rect 2763 13327 2805 13336
rect 1708 12452 1748 12461
rect 1611 12368 1653 12377
rect 1611 12328 1612 12368
rect 1652 12328 1653 12368
rect 1611 12319 1653 12328
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 1708 12209 1748 12412
rect 1900 12293 1940 12496
rect 2188 12491 2228 12500
rect 1996 12451 2188 12452
rect 2380 12487 2420 12496
rect 2476 13208 2516 13217
rect 1996 12412 2228 12451
rect 1899 12284 1941 12293
rect 1899 12244 1900 12284
rect 1940 12244 1941 12284
rect 1899 12235 1941 12244
rect 1996 12209 2036 12412
rect 2476 12377 2516 13168
rect 2571 12704 2613 12713
rect 2571 12664 2572 12704
rect 2612 12664 2613 12704
rect 2571 12655 2613 12664
rect 2572 12536 2612 12655
rect 2572 12487 2612 12496
rect 2668 12536 2708 12545
rect 2283 12368 2325 12377
rect 2380 12368 2420 12377
rect 2283 12328 2284 12368
rect 2324 12328 2380 12368
rect 2283 12319 2325 12328
rect 2380 12319 2420 12328
rect 2475 12368 2517 12377
rect 2475 12328 2476 12368
rect 2516 12328 2517 12368
rect 2475 12319 2517 12328
rect 2187 12284 2229 12293
rect 2187 12244 2188 12284
rect 2228 12244 2229 12284
rect 2187 12235 2229 12244
rect 1707 12200 1749 12209
rect 1707 12160 1708 12200
rect 1748 12160 1749 12200
rect 1707 12151 1749 12160
rect 1995 12200 2037 12209
rect 1995 12160 1996 12200
rect 2036 12160 2037 12200
rect 1995 12151 2037 12160
rect 1420 12076 1556 12116
rect 1419 11780 1461 11789
rect 1419 11740 1420 11780
rect 1460 11740 1461 11780
rect 1419 11731 1461 11740
rect 1420 11646 1460 11731
rect 1516 11192 1556 12076
rect 1804 11864 1844 11873
rect 2091 11864 2133 11873
rect 1844 11824 1940 11864
rect 1804 11815 1844 11824
rect 1228 11068 1364 11108
rect 1420 11152 1556 11192
rect 844 10940 884 10949
rect 844 10856 884 10900
rect 1132 10856 1172 10865
rect 844 10816 1132 10856
rect 1132 10807 1172 10816
rect 939 10352 981 10361
rect 939 10312 940 10352
rect 980 10312 981 10352
rect 939 10303 981 10312
rect 844 10268 884 10277
rect 844 9689 884 10228
rect 843 9680 885 9689
rect 843 9640 844 9680
rect 884 9640 885 9680
rect 843 9631 885 9640
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 844 8756 884 8765
rect 748 8716 844 8756
rect 844 8707 884 8716
rect 940 8588 980 10303
rect 1228 8756 1268 11068
rect 1324 10940 1364 10949
rect 1324 10445 1364 10900
rect 1323 10436 1365 10445
rect 1323 10396 1324 10436
rect 1364 10396 1365 10436
rect 1323 10387 1365 10396
rect 1420 9437 1460 11152
rect 1516 11024 1556 11033
rect 1900 11024 1940 11824
rect 2091 11824 2092 11864
rect 2132 11824 2133 11864
rect 2091 11815 2133 11824
rect 1995 11696 2037 11705
rect 1995 11656 1996 11696
rect 2036 11656 2037 11696
rect 1995 11647 2037 11656
rect 2092 11696 2132 11815
rect 1556 10984 1652 11024
rect 1516 10975 1556 10984
rect 1515 10352 1557 10361
rect 1515 10312 1516 10352
rect 1556 10312 1557 10352
rect 1515 10303 1557 10312
rect 1516 10218 1556 10303
rect 1612 10277 1652 10984
rect 1900 10975 1940 10984
rect 1996 10856 2036 11647
rect 1804 10816 2036 10856
rect 1611 10268 1653 10277
rect 1611 10228 1612 10268
rect 1652 10228 1653 10268
rect 1611 10219 1653 10228
rect 1708 10268 1748 10277
rect 1804 10268 1844 10816
rect 2092 10772 2132 11656
rect 1748 10228 1844 10268
rect 1996 10732 2132 10772
rect 2188 11696 2228 12235
rect 2668 11705 2708 12496
rect 1708 10219 1748 10228
rect 1515 9680 1557 9689
rect 1996 9680 2036 10732
rect 2188 10604 2228 11656
rect 2667 11696 2709 11705
rect 2667 11656 2668 11696
rect 2708 11656 2709 11696
rect 2667 11647 2709 11656
rect 2092 10564 2228 10604
rect 2284 11528 2324 11537
rect 2092 9848 2132 10564
rect 2188 10361 2228 10446
rect 2187 10352 2229 10361
rect 2187 10312 2188 10352
rect 2228 10312 2229 10352
rect 2187 10303 2229 10312
rect 2188 10184 2228 10193
rect 2284 10184 2324 11488
rect 2764 11024 2804 13327
rect 2860 12557 2900 13504
rect 2956 12713 2996 14008
rect 3051 14048 3093 14057
rect 3051 14008 3052 14048
rect 3092 14008 3093 14048
rect 3051 13999 3093 14008
rect 3052 13914 3092 13999
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3339 13376 3381 13385
rect 3339 13336 3340 13376
rect 3380 13336 3381 13376
rect 3339 13327 3381 13336
rect 3340 13208 3380 13327
rect 3340 13133 3380 13168
rect 3339 13124 3381 13133
rect 3339 13084 3340 13124
rect 3380 13084 3381 13124
rect 3339 13075 3381 13084
rect 3627 13040 3669 13049
rect 3627 13000 3628 13040
rect 3668 13000 3669 13040
rect 3627 12991 3669 13000
rect 2955 12704 2997 12713
rect 2955 12664 2956 12704
rect 2996 12664 2997 12704
rect 2955 12655 2997 12664
rect 2860 12517 2996 12557
rect 2859 12368 2901 12377
rect 2859 12328 2860 12368
rect 2900 12328 2901 12368
rect 2859 12319 2901 12328
rect 2860 12234 2900 12319
rect 2572 10984 2764 11024
rect 2475 10352 2517 10361
rect 2475 10312 2476 10352
rect 2516 10312 2517 10352
rect 2475 10303 2517 10312
rect 2228 10144 2324 10184
rect 2379 10184 2421 10193
rect 2379 10144 2380 10184
rect 2420 10144 2421 10184
rect 2188 10135 2228 10144
rect 2379 10135 2421 10144
rect 2476 10184 2516 10303
rect 2476 10135 2516 10144
rect 2380 10050 2420 10135
rect 2092 9808 2228 9848
rect 1515 9640 1516 9680
rect 1556 9640 1557 9680
rect 1515 9631 1557 9640
rect 1900 9640 2132 9680
rect 1516 9546 1556 9631
rect 1419 9428 1461 9437
rect 1419 9388 1420 9428
rect 1460 9388 1461 9428
rect 1419 9379 1461 9388
rect 1708 9428 1748 9437
rect 748 8548 980 8588
rect 1036 8716 1268 8756
rect 1324 9344 1364 9353
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 748 7244 788 8548
rect 844 7916 884 7925
rect 1036 7916 1076 8716
rect 1324 8672 1364 9304
rect 1708 8681 1748 9388
rect 1516 8672 1556 8681
rect 1324 8632 1516 8672
rect 1516 8623 1556 8632
rect 1707 8672 1749 8681
rect 1707 8632 1708 8672
rect 1748 8632 1749 8672
rect 1707 8623 1749 8632
rect 1132 8588 1172 8597
rect 1132 8177 1172 8548
rect 1227 8588 1269 8597
rect 1227 8548 1228 8588
rect 1268 8548 1269 8588
rect 1227 8539 1269 8548
rect 1131 8168 1173 8177
rect 1131 8128 1132 8168
rect 1172 8128 1173 8168
rect 1131 8119 1173 8128
rect 884 7876 1076 7916
rect 1228 7916 1268 8539
rect 1900 8168 1940 9640
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2092 9512 2132 9640
rect 2092 9463 2132 9472
rect 2188 9512 2228 9808
rect 1996 8765 2036 9463
rect 1995 8756 2037 8765
rect 1995 8716 1996 8756
rect 2036 8716 2037 8756
rect 1995 8707 2037 8716
rect 2188 8588 2228 9472
rect 844 7867 884 7876
rect 1228 7867 1268 7876
rect 1420 8128 1940 8168
rect 1036 7748 1076 7757
rect 940 7708 1036 7748
rect 844 7244 884 7253
rect 748 7204 844 7244
rect 844 7195 884 7204
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5144 692 5599
rect 844 5480 884 5489
rect 652 5095 692 5104
rect 748 5440 844 5480
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4304 692 4759
rect 652 4255 692 4264
rect 748 4220 788 5440
rect 844 5431 884 5440
rect 844 4892 884 4901
rect 940 4892 980 7708
rect 1036 7699 1076 7708
rect 1035 7580 1077 7589
rect 1035 7540 1036 7580
rect 1076 7540 1077 7580
rect 1035 7531 1077 7540
rect 1036 5732 1076 7531
rect 1036 5683 1076 5692
rect 1227 5564 1269 5573
rect 1227 5524 1228 5564
rect 1268 5524 1269 5564
rect 1227 5515 1269 5524
rect 1228 5430 1268 5515
rect 1420 5489 1460 8128
rect 1803 8000 1845 8009
rect 1803 7960 1804 8000
rect 1844 7960 1845 8000
rect 1803 7951 1845 7960
rect 1900 8000 1940 8128
rect 1900 7951 1940 7960
rect 1996 8548 2228 8588
rect 2284 9512 2324 9521
rect 1996 8000 2036 8548
rect 1612 7832 1652 7841
rect 1612 7160 1652 7792
rect 1804 7589 1844 7951
rect 1803 7580 1845 7589
rect 1803 7540 1804 7580
rect 1844 7540 1845 7580
rect 1803 7531 1845 7540
rect 1900 7160 1940 7169
rect 1612 7120 1900 7160
rect 1900 7111 1940 7120
rect 1516 7076 1556 7085
rect 1516 6665 1556 7036
rect 1996 6992 2036 7960
rect 1804 6952 2036 6992
rect 2092 8000 2132 8009
rect 1515 6656 1557 6665
rect 1515 6616 1516 6656
rect 1556 6616 1557 6656
rect 1515 6607 1557 6616
rect 1708 6320 1748 6329
rect 1515 5732 1557 5741
rect 1515 5692 1516 5732
rect 1556 5692 1557 5732
rect 1515 5683 1557 5692
rect 1419 5480 1461 5489
rect 1419 5440 1420 5480
rect 1460 5440 1461 5480
rect 1419 5431 1461 5440
rect 1516 4976 1556 5683
rect 1612 5648 1652 5657
rect 1708 5648 1748 6280
rect 1652 5608 1748 5648
rect 1612 5599 1652 5608
rect 1707 5480 1749 5489
rect 1707 5440 1708 5480
rect 1748 5440 1749 5480
rect 1707 5431 1749 5440
rect 1612 4976 1652 4985
rect 1516 4936 1612 4976
rect 884 4852 980 4892
rect 1420 4892 1460 4901
rect 1516 4892 1556 4936
rect 1612 4927 1652 4936
rect 1708 4976 1748 5431
rect 1460 4852 1556 4892
rect 844 4843 884 4852
rect 1420 4843 1460 4852
rect 1708 4808 1748 4936
rect 1612 4768 1748 4808
rect 1804 4976 1844 6952
rect 2092 6488 2132 7960
rect 2284 8000 2324 9472
rect 2380 8672 2420 8681
rect 2572 8672 2612 10984
rect 2764 10975 2804 10984
rect 2956 10856 2996 12517
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3435 11948 3477 11957
rect 3435 11908 3436 11948
rect 3476 11908 3477 11948
rect 3628 11948 3668 12991
rect 3820 11948 3860 15268
rect 3916 14309 3956 18115
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4780 17240 4820 18367
rect 4396 17200 4820 17240
rect 4203 16484 4245 16493
rect 4203 16444 4204 16484
rect 4244 16444 4245 16484
rect 4203 16435 4245 16444
rect 4011 16400 4053 16409
rect 4011 16360 4012 16400
rect 4052 16360 4053 16400
rect 4011 16351 4053 16360
rect 3915 14300 3957 14309
rect 3915 14260 3916 14300
rect 3956 14260 3957 14300
rect 3915 14251 3957 14260
rect 4012 14048 4052 16351
rect 4204 16350 4244 16435
rect 4396 16316 4436 17200
rect 5452 16997 5492 20728
rect 6123 20719 6165 20728
rect 5548 20600 5588 20609
rect 5548 20021 5588 20560
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 5547 20012 5589 20021
rect 5547 19972 5548 20012
rect 5588 19972 5589 20012
rect 5547 19963 5589 19972
rect 9003 20012 9045 20021
rect 9003 19972 9004 20012
rect 9044 19972 9045 20012
rect 9003 19963 9045 19972
rect 9004 19878 9044 19963
rect 9196 19844 9236 19853
rect 8812 19433 8852 19518
rect 6603 19424 6645 19433
rect 6603 19384 6604 19424
rect 6644 19384 6645 19424
rect 6603 19375 6645 19384
rect 7947 19424 7989 19433
rect 7947 19384 7948 19424
rect 7988 19384 7989 19424
rect 7947 19375 7989 19384
rect 8811 19424 8853 19433
rect 8811 19384 8812 19424
rect 8852 19384 8853 19424
rect 6604 19290 6644 19375
rect 7084 18584 7124 18593
rect 5932 18332 5972 18341
rect 5932 17669 5972 18292
rect 5931 17660 5973 17669
rect 5931 17620 5932 17660
rect 5972 17620 5973 17660
rect 5931 17611 5973 17620
rect 5451 16988 5493 16997
rect 5451 16948 5452 16988
rect 5492 16948 5493 16988
rect 5451 16939 5493 16948
rect 4875 16484 4917 16493
rect 4875 16444 4876 16484
rect 4916 16444 4917 16484
rect 4875 16435 4917 16444
rect 4396 16267 4436 16276
rect 4588 16148 4628 16157
rect 4628 16108 4820 16148
rect 4588 16099 4628 16108
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4299 15728 4341 15737
rect 4299 15688 4300 15728
rect 4340 15688 4341 15728
rect 4299 15679 4341 15688
rect 4396 15728 4436 15737
rect 4780 15728 4820 16108
rect 4436 15688 4820 15728
rect 4396 15679 4436 15688
rect 4203 15560 4245 15569
rect 4203 15520 4204 15560
rect 4244 15520 4245 15560
rect 4203 15511 4245 15520
rect 4300 15560 4340 15679
rect 4300 15511 4340 15520
rect 4492 15560 4532 15569
rect 4204 15426 4244 15511
rect 4492 15401 4532 15520
rect 4684 15560 4724 15571
rect 4684 15485 4724 15520
rect 4779 15560 4821 15569
rect 4779 15520 4780 15560
rect 4820 15520 4821 15560
rect 4779 15511 4821 15520
rect 4876 15560 4916 16435
rect 4683 15476 4725 15485
rect 4683 15436 4684 15476
rect 4724 15436 4725 15476
rect 4683 15427 4725 15436
rect 4780 15426 4820 15511
rect 4491 15392 4533 15401
rect 4491 15352 4492 15392
rect 4532 15352 4533 15392
rect 4491 15343 4533 15352
rect 4876 14720 4916 15520
rect 4972 16232 5012 16241
rect 4972 15392 5012 16192
rect 5835 16232 5877 16241
rect 5835 16192 5836 16232
rect 5876 16192 5877 16232
rect 5835 16183 5877 16192
rect 5836 16098 5876 16183
rect 5932 15980 5972 17611
rect 7084 16241 7124 18544
rect 7948 18584 7988 19375
rect 8524 19349 8564 19380
rect 8811 19375 8853 19384
rect 8523 19340 8565 19349
rect 8523 19300 8524 19340
rect 8564 19300 8565 19340
rect 8523 19291 8565 19300
rect 9003 19340 9045 19349
rect 9003 19300 9004 19340
rect 9044 19300 9045 19340
rect 9003 19291 9045 19300
rect 8332 19256 8372 19265
rect 8332 18929 8372 19216
rect 8524 19256 8564 19291
rect 8428 19088 8468 19097
rect 8331 18920 8373 18929
rect 8331 18880 8332 18920
rect 8372 18880 8373 18920
rect 8331 18871 8373 18880
rect 8332 18668 8372 18677
rect 8428 18668 8468 19048
rect 8524 18845 8564 19216
rect 8619 19256 8661 19265
rect 8619 19216 8620 19256
rect 8660 19216 8661 19256
rect 8619 19207 8661 19216
rect 8812 19256 8852 19265
rect 9004 19256 9044 19291
rect 9100 19265 9140 19350
rect 8852 19216 8948 19256
rect 8812 19207 8852 19216
rect 8620 19122 8660 19207
rect 8908 19004 8948 19216
rect 9004 19205 9044 19216
rect 9099 19256 9141 19265
rect 9099 19216 9100 19256
rect 9140 19216 9141 19256
rect 9099 19207 9141 19216
rect 8908 18964 9044 19004
rect 8811 18920 8853 18929
rect 8811 18880 8812 18920
rect 8852 18880 8853 18920
rect 8811 18871 8853 18880
rect 8523 18836 8565 18845
rect 8523 18796 8524 18836
rect 8564 18796 8565 18836
rect 8523 18787 8565 18796
rect 8372 18628 8468 18668
rect 8812 18668 8852 18871
rect 8907 18836 8949 18845
rect 8907 18796 8908 18836
rect 8948 18796 8949 18836
rect 8907 18787 8949 18796
rect 8332 18619 8372 18628
rect 8812 18619 8852 18628
rect 7948 18535 7988 18544
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 8523 18584 8565 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8716 18584 8756 18593
rect 8523 18535 8565 18544
rect 8620 18542 8660 18551
rect 7947 17828 7989 17837
rect 7947 17788 7948 17828
rect 7988 17788 7989 17828
rect 7947 17779 7989 17788
rect 7660 17744 7700 17753
rect 7660 16409 7700 17704
rect 7948 17744 7988 17779
rect 7948 17693 7988 17704
rect 8044 17669 8084 18535
rect 8524 18450 8564 18535
rect 8620 18173 8660 18502
rect 8619 18164 8661 18173
rect 8619 18124 8620 18164
rect 8660 18124 8661 18164
rect 8619 18115 8661 18124
rect 8619 17996 8661 18005
rect 8619 17956 8620 17996
rect 8660 17956 8661 17996
rect 8619 17947 8661 17956
rect 8332 17912 8372 17921
rect 8372 17872 8564 17912
rect 8332 17863 8372 17872
rect 8524 17744 8564 17872
rect 8620 17862 8660 17947
rect 8716 17912 8756 18544
rect 8908 18005 8948 18787
rect 9004 18752 9044 18964
rect 9004 18703 9044 18712
rect 9196 18677 9236 19804
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 21963 19592 22005 19601
rect 21963 19552 21964 19592
rect 22004 19552 22005 19592
rect 21963 19543 22005 19552
rect 11691 19508 11733 19517
rect 11691 19468 11692 19508
rect 11732 19468 11733 19508
rect 11691 19459 11733 19468
rect 9291 19424 9333 19433
rect 9291 19384 9292 19424
rect 9332 19384 9333 19424
rect 9291 19375 9333 19384
rect 9292 19256 9332 19375
rect 11692 19374 11732 19459
rect 21579 19340 21621 19349
rect 21579 19300 21580 19340
rect 21620 19300 21621 19340
rect 21579 19291 21621 19300
rect 21964 19340 22004 19543
rect 9292 19207 9332 19216
rect 9483 19256 9525 19265
rect 9483 19216 9484 19256
rect 9524 19216 9525 19256
rect 9483 19207 9525 19216
rect 9676 19256 9716 19265
rect 10539 19256 10581 19265
rect 9716 19216 9812 19256
rect 9676 19207 9716 19216
rect 9195 18668 9237 18677
rect 9195 18628 9196 18668
rect 9236 18628 9237 18668
rect 9195 18619 9237 18628
rect 9484 18668 9524 19207
rect 9484 18619 9524 18628
rect 9196 18500 9236 18619
rect 9196 18451 9236 18460
rect 9388 18584 9428 18593
rect 9004 18332 9044 18341
rect 8907 17996 8949 18005
rect 8907 17956 8908 17996
rect 8948 17956 8949 17996
rect 8907 17947 8949 17956
rect 8716 17872 8852 17912
rect 8524 17695 8564 17704
rect 8716 17744 8756 17753
rect 8043 17660 8085 17669
rect 8043 17620 8044 17660
rect 8084 17620 8085 17660
rect 8043 17611 8085 17620
rect 8044 17526 8084 17611
rect 7659 16400 7701 16409
rect 7659 16360 7660 16400
rect 7700 16360 7701 16400
rect 7659 16351 7701 16360
rect 6315 16232 6357 16241
rect 6315 16192 6316 16232
rect 6356 16192 6357 16232
rect 6315 16183 6357 16192
rect 7083 16232 7125 16241
rect 7083 16192 7084 16232
rect 7124 16192 7125 16232
rect 7083 16183 7125 16192
rect 5836 15940 5972 15980
rect 5068 15392 5108 15401
rect 4972 15352 5068 15392
rect 5068 15343 5108 15352
rect 5068 14720 5108 14729
rect 4876 14680 5068 14720
rect 4779 14636 4821 14645
rect 4779 14596 4780 14636
rect 4820 14596 4821 14636
rect 4779 14587 4821 14596
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4299 14132 4341 14141
rect 4299 14092 4300 14132
rect 4340 14092 4341 14132
rect 4299 14083 4341 14092
rect 3628 11908 3669 11948
rect 3435 11899 3477 11908
rect 3339 11864 3381 11873
rect 3339 11824 3340 11864
rect 3380 11824 3381 11864
rect 3339 11815 3381 11824
rect 3340 11696 3380 11815
rect 3340 11647 3380 11656
rect 3436 11453 3476 11899
rect 3531 11864 3573 11873
rect 3531 11824 3532 11864
rect 3572 11824 3573 11864
rect 3531 11815 3573 11824
rect 3435 11444 3477 11453
rect 3435 11404 3436 11444
rect 3476 11404 3477 11444
rect 3435 11395 3477 11404
rect 2764 10816 2996 10856
rect 2668 10361 2708 10446
rect 2667 10352 2709 10361
rect 2667 10312 2668 10352
rect 2708 10312 2709 10352
rect 2667 10303 2709 10312
rect 2420 8632 2612 8672
rect 2668 10184 2708 10193
rect 2764 10184 2804 10816
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3435 10436 3477 10445
rect 3435 10396 3436 10436
rect 3476 10396 3477 10436
rect 3435 10387 3477 10396
rect 3148 10352 3188 10361
rect 2708 10144 2804 10184
rect 2956 10184 2996 10193
rect 2380 8623 2420 8632
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 2379 8168 2421 8177
rect 2379 8128 2380 8168
rect 2420 8128 2421 8168
rect 2379 8119 2421 8128
rect 2380 8034 2420 8119
rect 2284 7951 2324 7960
rect 2476 8000 2516 8455
rect 2476 7951 2516 7960
rect 2572 8000 2612 8009
rect 2572 7841 2612 7960
rect 2668 8000 2708 10144
rect 2860 10142 2900 10151
rect 2859 10102 2860 10109
rect 2900 10102 2901 10109
rect 2859 10100 2901 10102
rect 2859 10060 2860 10100
rect 2900 10060 2901 10100
rect 2859 10051 2901 10060
rect 2860 10007 2900 10051
rect 2859 9680 2901 9689
rect 2859 9640 2860 9680
rect 2900 9640 2901 9680
rect 2859 9631 2901 9640
rect 2860 9527 2900 9631
rect 2956 9521 2996 10144
rect 3148 10109 3188 10312
rect 3339 10268 3381 10277
rect 3339 10228 3340 10268
rect 3380 10228 3381 10268
rect 3339 10219 3381 10228
rect 3340 10134 3380 10219
rect 3147 10100 3189 10109
rect 3052 10060 3148 10100
rect 3188 10060 3189 10100
rect 2860 9344 2900 9487
rect 2955 9512 2997 9521
rect 2955 9472 2956 9512
rect 2996 9472 2997 9512
rect 2955 9463 2997 9472
rect 2764 9304 2900 9344
rect 2764 8849 2804 9304
rect 3052 9260 3092 10060
rect 3147 10051 3189 10060
rect 3148 9512 3188 9523
rect 3148 9437 3188 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3147 9428 3189 9437
rect 3147 9388 3148 9428
rect 3188 9388 3189 9428
rect 3147 9379 3189 9388
rect 3244 9378 3284 9463
rect 3436 9269 3476 10387
rect 3532 9689 3572 11815
rect 3629 11780 3669 11908
rect 3819 11908 3860 11948
rect 3916 14008 4012 14048
rect 3819 11864 3859 11908
rect 3916 11873 3956 14008
rect 4012 13999 4052 14008
rect 4300 14048 4340 14083
rect 4300 13973 4340 14008
rect 4395 14048 4437 14057
rect 4395 14008 4396 14048
rect 4436 14008 4437 14048
rect 4395 13999 4437 14008
rect 4299 13964 4341 13973
rect 4299 13924 4300 13964
rect 4340 13924 4341 13964
rect 4299 13915 4341 13924
rect 4300 13884 4340 13915
rect 4396 13460 4436 13999
rect 4683 13796 4725 13805
rect 4683 13756 4684 13796
rect 4724 13756 4725 13796
rect 4683 13747 4725 13756
rect 4684 13662 4724 13747
rect 4492 13460 4532 13469
rect 4396 13420 4492 13460
rect 4492 13411 4532 13420
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4587 12704 4629 12713
rect 4587 12664 4588 12704
rect 4628 12664 4629 12704
rect 4587 12655 4629 12664
rect 4588 12570 4628 12655
rect 4491 12536 4533 12545
rect 4491 12496 4492 12536
rect 4532 12496 4533 12536
rect 4491 12487 4533 12496
rect 4684 12536 4724 12545
rect 3915 11864 3957 11873
rect 3819 11824 3860 11864
rect 3628 11740 3669 11780
rect 3628 11696 3668 11740
rect 3628 11621 3668 11656
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 3627 11612 3669 11621
rect 3627 11572 3628 11612
rect 3668 11572 3669 11612
rect 3627 11563 3669 11572
rect 3724 11562 3764 11647
rect 3627 11444 3669 11453
rect 3627 11404 3628 11444
rect 3668 11404 3669 11444
rect 3627 11395 3669 11404
rect 3531 9680 3573 9689
rect 3531 9640 3532 9680
rect 3572 9640 3573 9680
rect 3531 9631 3573 9640
rect 3628 9605 3668 11395
rect 3820 11117 3860 11824
rect 3915 11824 3916 11864
rect 3956 11824 3957 11864
rect 3915 11815 3957 11824
rect 4012 11864 4052 11873
rect 4052 11824 4148 11864
rect 4012 11815 4052 11824
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 3916 11192 3956 11647
rect 3916 11143 3956 11152
rect 3819 11108 3861 11117
rect 3819 11068 3820 11108
rect 3860 11068 3861 11108
rect 3819 11059 3861 11068
rect 3627 9596 3669 9605
rect 3627 9556 3628 9596
rect 3668 9556 3669 9596
rect 3627 9547 3669 9556
rect 3724 9512 3764 9521
rect 3820 9512 3860 11059
rect 4108 11024 4148 11824
rect 4492 11696 4532 12487
rect 4684 12368 4724 12496
rect 4780 12536 4820 14587
rect 4876 14477 4916 14680
rect 5068 14671 5108 14680
rect 5259 14720 5301 14729
rect 5259 14680 5260 14720
rect 5300 14680 5301 14720
rect 5259 14671 5301 14680
rect 5163 14636 5205 14645
rect 5163 14596 5164 14636
rect 5204 14596 5205 14636
rect 5163 14587 5205 14596
rect 5164 14502 5204 14587
rect 4875 14468 4917 14477
rect 4875 14428 4876 14468
rect 4916 14428 4917 14468
rect 4875 14419 4917 14428
rect 5260 14141 5300 14671
rect 5259 14132 5301 14141
rect 5259 14092 5260 14132
rect 5300 14092 5301 14132
rect 5259 14083 5301 14092
rect 5068 14048 5108 14057
rect 4875 13292 4917 13301
rect 4875 13252 4876 13292
rect 4916 13252 4917 13292
rect 4875 13243 4917 13252
rect 4780 12487 4820 12496
rect 4876 12368 4916 13243
rect 5068 12713 5108 14008
rect 5452 14048 5492 14057
rect 5452 13385 5492 14008
rect 5356 13376 5396 13385
rect 5163 13208 5205 13217
rect 5163 13168 5164 13208
rect 5204 13168 5205 13208
rect 5163 13159 5205 13168
rect 5067 12704 5109 12713
rect 5067 12664 5068 12704
rect 5108 12664 5109 12704
rect 5067 12655 5109 12664
rect 4684 12328 4916 12368
rect 4492 11647 4532 11656
rect 4588 11824 5012 11864
rect 4588 11612 4628 11824
rect 4588 11563 4628 11572
rect 4684 11696 4724 11705
rect 4684 11537 4724 11656
rect 4780 11696 4820 11705
rect 4203 11528 4245 11537
rect 4203 11488 4204 11528
rect 4244 11488 4245 11528
rect 4203 11479 4245 11488
rect 4683 11528 4725 11537
rect 4683 11488 4684 11528
rect 4724 11488 4725 11528
rect 4683 11479 4725 11488
rect 4108 10975 4148 10984
rect 4204 10772 4244 11479
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4780 11360 4820 11656
rect 4972 11696 5012 11824
rect 4972 11647 5012 11656
rect 5067 11612 5109 11621
rect 5067 11572 5068 11612
rect 5108 11572 5109 11612
rect 5067 11563 5109 11572
rect 4780 11320 5012 11360
rect 4352 11311 4720 11320
rect 4587 11192 4629 11201
rect 4587 11152 4588 11192
rect 4628 11152 4629 11192
rect 4587 11143 4629 11152
rect 4299 11108 4341 11117
rect 4299 11068 4300 11108
rect 4340 11068 4341 11108
rect 4299 11059 4341 11068
rect 4300 11024 4340 11059
rect 4300 10973 4340 10984
rect 4204 10193 4244 10732
rect 4203 10184 4245 10193
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 4588 10025 4628 11143
rect 4972 11108 5012 11320
rect 4972 11059 5012 11068
rect 4875 11024 4917 11033
rect 4875 10984 4876 11024
rect 4916 10984 4917 11024
rect 4875 10975 4917 10984
rect 5068 11024 5108 11563
rect 5068 10975 5108 10984
rect 4876 10277 4916 10975
rect 5067 10352 5109 10361
rect 5067 10312 5068 10352
rect 5108 10312 5109 10352
rect 5067 10303 5109 10312
rect 4875 10268 4917 10277
rect 4875 10228 4876 10268
rect 4916 10228 4917 10268
rect 4875 10219 4917 10228
rect 4876 10100 4916 10219
rect 4876 10060 5012 10100
rect 4587 10016 4629 10025
rect 4587 9976 4588 10016
rect 4628 9976 4629 10016
rect 4587 9967 4629 9976
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4492 9605 4532 9690
rect 4491 9596 4533 9605
rect 4491 9556 4492 9596
rect 4532 9556 4533 9596
rect 4491 9547 4533 9556
rect 4779 9596 4821 9605
rect 4779 9556 4780 9596
rect 4820 9556 4821 9596
rect 4779 9547 4821 9556
rect 3916 9512 3956 9521
rect 4299 9512 4341 9521
rect 3820 9472 3916 9512
rect 3956 9472 4244 9512
rect 3724 9428 3764 9472
rect 3916 9463 3956 9472
rect 3532 9388 3764 9428
rect 3532 9386 3572 9388
rect 3532 9337 3572 9346
rect 2956 9220 3092 9260
rect 3435 9260 3477 9269
rect 3435 9220 3436 9260
rect 3476 9220 3477 9260
rect 2763 8840 2805 8849
rect 2763 8800 2764 8840
rect 2804 8800 2805 8840
rect 2763 8791 2805 8800
rect 2764 8000 2804 8009
rect 2668 7960 2764 8000
rect 2571 7832 2613 7841
rect 2571 7792 2572 7832
rect 2612 7792 2613 7832
rect 2571 7783 2613 7792
rect 2668 7328 2708 7960
rect 2764 7951 2804 7960
rect 2956 8000 2996 9220
rect 3435 9211 3477 9220
rect 3627 9260 3669 9269
rect 3627 9220 3628 9260
rect 3668 9220 3669 9260
rect 3627 9211 3669 9220
rect 3820 9260 3860 9269
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3435 8840 3477 8849
rect 3435 8800 3436 8840
rect 3476 8800 3477 8840
rect 3435 8791 3477 8800
rect 2763 7832 2805 7841
rect 2763 7792 2764 7832
rect 2804 7792 2805 7832
rect 2763 7783 2805 7792
rect 2764 7698 2804 7783
rect 2572 7288 2708 7328
rect 2283 7076 2325 7085
rect 2283 7036 2284 7076
rect 2324 7036 2325 7076
rect 2283 7027 2325 7036
rect 2187 6656 2229 6665
rect 2187 6616 2188 6656
rect 2228 6616 2229 6656
rect 2187 6607 2229 6616
rect 2188 6522 2228 6607
rect 2092 6439 2132 6448
rect 2284 6488 2324 7027
rect 2284 6439 2324 6448
rect 2380 6488 2420 6497
rect 2572 6488 2612 7288
rect 2956 7169 2996 7960
rect 3051 8000 3093 8009
rect 3051 7960 3052 8000
rect 3092 7960 3093 8000
rect 3051 7951 3093 7960
rect 3436 8000 3476 8791
rect 3531 8756 3573 8765
rect 3531 8716 3532 8756
rect 3572 8716 3573 8756
rect 3531 8707 3573 8716
rect 3532 8622 3572 8707
rect 3476 7960 3572 8000
rect 3436 7951 3476 7960
rect 3052 7866 3092 7951
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 2764 7160 2804 7169
rect 2380 6329 2420 6448
rect 2476 6448 2572 6488
rect 2379 6320 2421 6329
rect 2379 6280 2380 6320
rect 2420 6280 2421 6320
rect 2379 6271 2421 6280
rect 2476 6152 2516 6448
rect 2572 6439 2612 6448
rect 2668 7120 2764 7160
rect 2571 6320 2613 6329
rect 2571 6280 2572 6320
rect 2612 6280 2613 6320
rect 2571 6271 2613 6280
rect 2572 6186 2612 6271
rect 2380 6112 2516 6152
rect 2187 5564 2229 5573
rect 2187 5524 2188 5564
rect 2228 5524 2229 5564
rect 2187 5515 2229 5524
rect 2188 5144 2228 5515
rect 2188 5095 2228 5104
rect 2283 5144 2325 5153
rect 2283 5104 2284 5144
rect 2324 5104 2325 5144
rect 2380 5144 2420 6112
rect 2476 5648 2516 5657
rect 2668 5648 2708 7120
rect 2764 7111 2804 7120
rect 2955 7160 2997 7169
rect 2955 7120 2956 7160
rect 2996 7120 2997 7160
rect 2955 7111 2997 7120
rect 2956 6656 2996 7111
rect 2764 6616 2996 6656
rect 2764 6488 2804 6616
rect 3532 6497 3572 7960
rect 3628 6581 3668 9211
rect 3820 8513 3860 9220
rect 3819 8504 3861 8513
rect 3819 8464 3820 8504
rect 3860 8464 3861 8504
rect 3819 8455 3861 8464
rect 3724 8000 3764 8009
rect 3724 7757 3764 7960
rect 3819 8000 3861 8009
rect 3819 7960 3820 8000
rect 3860 7960 3956 8000
rect 3819 7951 3861 7960
rect 3820 7866 3860 7951
rect 3723 7748 3765 7757
rect 3723 7708 3724 7748
rect 3764 7708 3765 7748
rect 3723 7699 3765 7708
rect 3916 7412 3956 7960
rect 4204 7916 4244 9472
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4396 9512 4436 9521
rect 4300 9378 4340 9463
rect 4396 8513 4436 9472
rect 4588 9512 4628 9521
rect 4491 9428 4533 9437
rect 4491 9388 4492 9428
rect 4532 9388 4533 9428
rect 4491 9379 4533 9388
rect 4492 8681 4532 9379
rect 4588 9353 4628 9472
rect 4780 9462 4820 9547
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 4587 9344 4629 9353
rect 4587 9304 4588 9344
rect 4628 9304 4629 9344
rect 4587 9295 4629 9304
rect 4779 8840 4821 8849
rect 4779 8800 4780 8840
rect 4820 8800 4821 8840
rect 4779 8791 4821 8800
rect 4491 8672 4533 8681
rect 4491 8632 4492 8672
rect 4532 8632 4533 8672
rect 4491 8623 4533 8632
rect 4780 8672 4820 8791
rect 4780 8623 4820 8632
rect 4876 8588 4916 9463
rect 4972 8849 5012 10060
rect 5068 9512 5108 10303
rect 5164 9680 5204 13159
rect 5356 13133 5396 13336
rect 5451 13376 5493 13385
rect 5451 13336 5452 13376
rect 5492 13336 5493 13376
rect 5451 13327 5493 13336
rect 5355 13124 5397 13133
rect 5355 13084 5356 13124
rect 5396 13084 5397 13124
rect 5355 13075 5397 13084
rect 5356 12536 5396 13075
rect 5356 12487 5396 12496
rect 5355 12368 5397 12377
rect 5355 12328 5356 12368
rect 5396 12328 5397 12368
rect 5355 12319 5397 12328
rect 5356 11696 5396 12319
rect 5356 11647 5396 11656
rect 5259 10352 5301 10361
rect 5259 10312 5260 10352
rect 5300 10312 5301 10352
rect 5259 10303 5301 10312
rect 5260 10218 5300 10303
rect 5164 9640 5300 9680
rect 5164 9512 5204 9521
rect 5068 9472 5164 9512
rect 5164 9463 5204 9472
rect 4971 8840 5013 8849
rect 4971 8800 4972 8840
rect 5012 8800 5013 8840
rect 4971 8791 5013 8800
rect 4971 8672 5013 8681
rect 4971 8632 4972 8672
rect 5012 8632 5013 8672
rect 4971 8623 5013 8632
rect 4876 8539 4916 8548
rect 4972 8538 5012 8623
rect 4395 8504 4437 8513
rect 4395 8464 4396 8504
rect 4436 8464 4437 8504
rect 4395 8455 4437 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4684 8168 4724 8177
rect 4724 8128 5108 8168
rect 4684 8119 4724 8128
rect 5068 8084 5108 8128
rect 5068 8035 5108 8044
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4780 8000 4820 8009
rect 3916 7363 3956 7372
rect 4012 7876 4244 7916
rect 3627 6572 3669 6581
rect 3627 6532 3628 6572
rect 3668 6532 3669 6572
rect 3627 6523 3669 6532
rect 3915 6572 3957 6581
rect 3915 6532 3916 6572
rect 3956 6532 3957 6572
rect 3915 6523 3957 6532
rect 3531 6488 3573 6497
rect 2764 6439 2804 6448
rect 2870 6469 2910 6478
rect 3531 6448 3532 6488
rect 3572 6448 3573 6488
rect 3531 6439 3573 6448
rect 2870 6068 2910 6429
rect 3112 6068 3480 6077
rect 2870 6028 2996 6068
rect 2956 5741 2996 6028
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 2955 5732 2997 5741
rect 2955 5692 2956 5732
rect 2996 5692 2997 5732
rect 2955 5683 2997 5692
rect 2516 5608 2804 5648
rect 2476 5599 2516 5608
rect 2380 5104 2516 5144
rect 2283 5095 2325 5104
rect 1804 4808 1844 4936
rect 1900 4976 1940 4985
rect 2092 4976 2132 4985
rect 1940 4936 2092 4976
rect 1900 4927 1940 4936
rect 2092 4927 2132 4936
rect 2284 4976 2324 5095
rect 2284 4927 2324 4936
rect 2380 4976 2420 4985
rect 1804 4768 1940 4808
rect 1228 4724 1268 4733
rect 844 4220 884 4229
rect 748 4180 844 4220
rect 844 4171 884 4180
rect 1228 4220 1268 4684
rect 1228 4171 1268 4180
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 1036 3834 1076 3919
rect 1323 3548 1365 3557
rect 1323 3508 1324 3548
rect 1364 3508 1365 3548
rect 1323 3499 1365 3508
rect 1324 3414 1364 3499
rect 1131 3380 1173 3389
rect 1131 3340 1132 3380
rect 1172 3340 1173 3380
rect 1131 3331 1173 3340
rect 1132 3246 1172 3331
rect 1612 3221 1652 4768
rect 1804 4304 1844 4313
rect 1708 4264 1804 4304
rect 1708 3464 1748 4264
rect 1804 4255 1844 4264
rect 1708 3415 1748 3424
rect 1900 3305 1940 4768
rect 2380 4388 2420 4936
rect 2380 4339 2420 4348
rect 2380 4136 2420 4145
rect 2476 4136 2516 5104
rect 2764 5069 2804 5608
rect 3532 5480 3572 6439
rect 3820 6236 3860 6245
rect 3724 6196 3820 6236
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 3628 5598 3668 5683
rect 3340 5440 3572 5480
rect 2763 5060 2805 5069
rect 2763 5020 2764 5060
rect 2804 5020 2805 5060
rect 2763 5011 2805 5020
rect 2420 4096 2516 4136
rect 2572 4136 2612 4145
rect 1899 3296 1941 3305
rect 1899 3256 1900 3296
rect 1940 3256 1941 3296
rect 1899 3247 1941 3256
rect 940 3212 980 3221
rect 651 3128 693 3137
rect 651 3088 652 3128
rect 692 3088 693 3128
rect 651 3079 693 3088
rect 652 2876 692 3079
rect 652 2827 692 2836
rect 844 2708 884 2717
rect 940 2708 980 3172
rect 1611 3212 1653 3221
rect 1611 3172 1612 3212
rect 1652 3172 1653 3212
rect 1611 3163 1653 3172
rect 1516 2792 1556 2801
rect 884 2668 980 2708
rect 1228 2752 1516 2792
rect 1228 2708 1268 2752
rect 1516 2743 1556 2752
rect 844 2659 884 2668
rect 1228 2659 1268 2668
rect 1707 2708 1749 2717
rect 1707 2668 1708 2708
rect 1748 2668 1749 2708
rect 1707 2659 1749 2668
rect 1708 2574 1748 2659
rect 2380 2633 2420 4096
rect 2572 3977 2612 4096
rect 2668 4136 2708 4145
rect 2668 4061 2708 4096
rect 2667 4052 2709 4061
rect 2667 4012 2668 4052
rect 2708 4012 2709 4052
rect 2667 4003 2709 4012
rect 2571 3968 2613 3977
rect 2571 3928 2572 3968
rect 2612 3928 2613 3968
rect 2571 3919 2613 3928
rect 2668 3632 2708 4003
rect 2476 3592 2708 3632
rect 2476 3389 2516 3592
rect 2572 3464 2612 3473
rect 2764 3464 2804 5011
rect 3340 4808 3380 5440
rect 3435 5312 3477 5321
rect 3435 5272 3436 5312
rect 3476 5272 3477 5312
rect 3435 5263 3477 5272
rect 3436 4985 3476 5263
rect 3531 5228 3573 5237
rect 3531 5188 3532 5228
rect 3572 5188 3573 5228
rect 3531 5179 3573 5188
rect 3532 5060 3572 5179
rect 3532 5011 3572 5020
rect 3435 4976 3477 4985
rect 3435 4936 3436 4976
rect 3476 4936 3477 4976
rect 3435 4927 3477 4936
rect 3628 4976 3668 4985
rect 3724 4976 3764 6196
rect 3820 6187 3860 6196
rect 3916 5480 3956 6523
rect 3668 4936 3764 4976
rect 3820 5440 3956 5480
rect 3820 4976 3860 5440
rect 4012 5321 4052 7876
rect 4108 7748 4148 7757
rect 4108 7160 4148 7708
rect 4204 7328 4244 7876
rect 4588 7866 4628 7951
rect 4204 7288 4436 7328
rect 4204 7160 4244 7169
rect 4108 7120 4204 7160
rect 4204 7111 4244 7120
rect 4300 7085 4340 7170
rect 4396 7160 4436 7288
rect 4396 7111 4436 7120
rect 4780 7085 4820 7960
rect 4876 8000 4916 8009
rect 4876 7412 4916 7960
rect 5163 7748 5205 7757
rect 5163 7708 5164 7748
rect 5204 7708 5205 7748
rect 5163 7699 5205 7708
rect 5068 7412 5108 7421
rect 4876 7372 5068 7412
rect 5068 7363 5108 7372
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4971 7111 5013 7120
rect 5164 7160 5204 7699
rect 5164 7111 5204 7120
rect 4299 7076 4341 7085
rect 4299 7036 4300 7076
rect 4340 7036 4341 7076
rect 4299 7027 4341 7036
rect 4779 7076 4821 7085
rect 4779 7036 4780 7076
rect 4820 7036 4821 7076
rect 4779 7027 4821 7036
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 4203 6572 4245 6581
rect 4203 6532 4204 6572
rect 4244 6532 4245 6572
rect 4203 6523 4245 6532
rect 4108 6488 4148 6497
rect 4108 5741 4148 6448
rect 4204 6488 4244 6523
rect 4204 6437 4244 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 4492 6354 4532 6439
rect 4972 6077 5012 7111
rect 5068 6488 5108 6497
rect 4203 6068 4245 6077
rect 4203 6028 4204 6068
rect 4244 6028 4245 6068
rect 4203 6019 4245 6028
rect 4971 6068 5013 6077
rect 4971 6028 4972 6068
rect 5012 6028 5013 6068
rect 4971 6019 5013 6028
rect 4107 5732 4149 5741
rect 4107 5692 4108 5732
rect 4148 5692 4149 5732
rect 4107 5683 4149 5692
rect 4011 5312 4053 5321
rect 4011 5272 4012 5312
rect 4052 5272 4053 5312
rect 4011 5263 4053 5272
rect 3915 5144 3957 5153
rect 4204 5144 4244 6019
rect 5068 5909 5108 6448
rect 5067 5900 5109 5909
rect 5067 5860 5068 5900
rect 5108 5860 5109 5900
rect 5067 5851 5109 5860
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3915 5104 3916 5144
rect 3956 5104 3957 5144
rect 3915 5095 3957 5104
rect 4012 5104 4244 5144
rect 3916 5060 3956 5095
rect 3916 5009 3956 5020
rect 3628 4927 3668 4936
rect 3820 4927 3860 4936
rect 4012 4976 4052 5104
rect 4299 5060 4341 5069
rect 4299 5020 4300 5060
rect 4340 5020 4341 5060
rect 4299 5011 4341 5020
rect 3340 4768 3572 4808
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 3051 4136 3093 4145
rect 2612 3424 2804 3464
rect 2860 4094 2900 4103
rect 3051 4096 3052 4136
rect 3092 4096 3093 4136
rect 3051 4087 3093 4096
rect 3148 4136 3188 4145
rect 2572 3415 2612 3424
rect 2475 3380 2517 3389
rect 2860 3380 2900 4054
rect 3052 4002 3092 4087
rect 2956 3968 2996 3977
rect 2956 3557 2996 3928
rect 2955 3548 2997 3557
rect 2955 3508 2956 3548
rect 2996 3508 2997 3548
rect 2955 3499 2997 3508
rect 3148 3380 3188 4096
rect 3532 4136 3572 4768
rect 3819 4304 3861 4313
rect 3819 4264 3820 4304
rect 3860 4264 3861 4304
rect 3819 4255 3861 4264
rect 3532 4087 3572 4096
rect 3820 4136 3860 4255
rect 3820 4087 3860 4096
rect 3723 4052 3765 4061
rect 3723 4012 3724 4052
rect 3764 4012 3765 4052
rect 3723 4003 3765 4012
rect 3915 4052 3957 4061
rect 3915 4012 3916 4052
rect 3956 4012 3957 4052
rect 3915 4003 3957 4012
rect 3531 3968 3573 3977
rect 3531 3928 3532 3968
rect 3572 3928 3573 3968
rect 3531 3919 3573 3928
rect 2475 3340 2476 3380
rect 2516 3340 2517 3380
rect 2475 3331 2517 3340
rect 2764 3340 2900 3380
rect 2956 3340 3188 3380
rect 2379 2624 2421 2633
rect 2379 2584 2380 2624
rect 2420 2584 2421 2624
rect 2379 2575 2421 2584
rect 2476 2624 2516 3331
rect 2667 3296 2709 3305
rect 2667 3256 2668 3296
rect 2708 3256 2709 3296
rect 2667 3247 2709 3256
rect 2571 3212 2613 3221
rect 2571 3172 2572 3212
rect 2612 3172 2613 3212
rect 2571 3163 2613 3172
rect 2476 2575 2516 2584
rect 2572 2624 2612 3163
rect 2572 2575 2612 2584
rect 2668 2624 2708 3247
rect 2764 2900 2804 3340
rect 2764 2860 2900 2900
rect 2668 2575 2708 2584
rect 2764 2624 2804 2633
rect 2860 2624 2900 2860
rect 2956 2876 2996 3340
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 3052 2876 3092 2885
rect 3532 2876 3572 3919
rect 3724 3632 3764 4003
rect 3916 3918 3956 4003
rect 4012 3977 4052 4936
rect 4300 4926 4340 5011
rect 4683 4976 4725 4985
rect 4683 4936 4684 4976
rect 4724 4936 4725 4976
rect 4683 4927 4725 4936
rect 5164 4976 5204 4985
rect 5260 4976 5300 9640
rect 5452 8000 5492 8009
rect 5452 7328 5492 7960
rect 5548 7328 5588 7337
rect 5452 7288 5548 7328
rect 5548 7279 5588 7288
rect 5204 4936 5300 4976
rect 5452 6488 5492 6497
rect 5164 4927 5204 4936
rect 4204 4304 4244 4313
rect 4011 3968 4053 3977
rect 4011 3928 4012 3968
rect 4052 3928 4053 3968
rect 4011 3919 4053 3928
rect 3724 3583 3764 3592
rect 4204 3464 4244 4264
rect 4395 4304 4437 4313
rect 4395 4264 4396 4304
rect 4436 4264 4437 4304
rect 4395 4255 4437 4264
rect 4396 4136 4436 4255
rect 4491 4220 4533 4229
rect 4491 4180 4492 4220
rect 4532 4180 4533 4220
rect 4491 4171 4533 4180
rect 4396 4087 4436 4096
rect 4492 4086 4532 4171
rect 4588 4136 4628 4145
rect 4588 3977 4628 4096
rect 4587 3968 4629 3977
rect 4587 3928 4588 3968
rect 4628 3928 4629 3968
rect 4684 3968 4724 4927
rect 5452 4808 5492 6448
rect 5739 5648 5781 5657
rect 5739 5608 5740 5648
rect 5780 5608 5781 5648
rect 5739 5599 5781 5608
rect 5740 5069 5780 5599
rect 5739 5060 5781 5069
rect 5739 5020 5740 5060
rect 5780 5020 5781 5060
rect 5739 5011 5781 5020
rect 5836 4976 5876 15940
rect 6316 14048 6356 16183
rect 6795 16064 6837 16073
rect 6795 16024 6796 16064
rect 6836 16024 6837 16064
rect 6795 16015 6837 16024
rect 6987 16064 7029 16073
rect 6987 16024 6988 16064
rect 7028 16024 7029 16064
rect 6987 16015 7029 16024
rect 6796 15905 6836 16015
rect 6795 15896 6837 15905
rect 6795 15856 6796 15896
rect 6836 15856 6837 15896
rect 6795 15847 6837 15856
rect 6219 13376 6261 13385
rect 6219 13336 6220 13376
rect 6260 13336 6261 13376
rect 6219 13327 6261 13336
rect 6220 13242 6260 13327
rect 6028 13208 6068 13217
rect 6028 12980 6068 13168
rect 6316 12980 6356 14008
rect 6603 13796 6645 13805
rect 6603 13756 6604 13796
rect 6644 13756 6645 13796
rect 6603 13747 6645 13756
rect 6604 13208 6644 13747
rect 6699 13292 6741 13301
rect 6699 13252 6700 13292
rect 6740 13252 6741 13292
rect 6699 13243 6741 13252
rect 6604 13159 6644 13168
rect 6700 13158 6740 13243
rect 6796 13208 6836 15847
rect 6988 15485 7028 16015
rect 8716 15905 8756 17704
rect 8812 17249 8852 17872
rect 8811 17240 8853 17249
rect 8811 17200 8812 17240
rect 8852 17200 8853 17240
rect 8811 17191 8853 17200
rect 8715 15896 8757 15905
rect 8715 15856 8716 15896
rect 8756 15856 8757 15896
rect 8715 15847 8757 15856
rect 6987 15476 7029 15485
rect 6987 15436 6988 15476
rect 7028 15436 7029 15476
rect 6987 15427 7029 15436
rect 9004 15401 9044 18292
rect 9388 16493 9428 18544
rect 9579 18584 9621 18593
rect 9579 18544 9580 18584
rect 9620 18544 9621 18584
rect 9579 18535 9621 18544
rect 9580 17837 9620 18535
rect 9772 18416 9812 19216
rect 10539 19216 10540 19256
rect 10580 19216 10581 19256
rect 10539 19207 10581 19216
rect 10540 19122 10580 19207
rect 11692 19088 11732 19097
rect 11692 18593 11732 19048
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 11691 18584 11733 18593
rect 11691 18544 11692 18584
rect 11732 18544 11733 18584
rect 11691 18535 11733 18544
rect 9772 18367 9812 18376
rect 21484 18500 21524 18509
rect 21484 18257 21524 18460
rect 21483 18248 21525 18257
rect 21483 18208 21484 18248
rect 21524 18208 21525 18248
rect 21483 18199 21525 18208
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 9579 17828 9621 17837
rect 9579 17788 9580 17828
rect 9620 17788 9621 17828
rect 9579 17779 9621 17788
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 9387 16484 9429 16493
rect 9387 16444 9388 16484
rect 9428 16444 9429 16484
rect 9387 16435 9429 16444
rect 21580 15989 21620 19291
rect 21771 19088 21813 19097
rect 21771 19048 21772 19088
rect 21812 19048 21813 19088
rect 21771 19039 21813 19048
rect 21772 18954 21812 19039
rect 21676 18332 21716 18341
rect 21676 17753 21716 18292
rect 21868 18332 21908 18343
rect 21868 18257 21908 18292
rect 21867 18248 21909 18257
rect 21867 18208 21868 18248
rect 21908 18208 21909 18248
rect 21867 18199 21909 18208
rect 21675 17744 21717 17753
rect 21675 17704 21676 17744
rect 21716 17704 21717 17744
rect 21675 17695 21717 17704
rect 21964 16157 22004 19300
rect 22060 18677 22100 22987
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 28012 22364 28052 22373
rect 28012 22205 28052 22324
rect 27531 22196 27573 22205
rect 27531 22156 27532 22196
rect 27572 22156 27573 22196
rect 27531 22147 27573 22156
rect 28011 22196 28053 22205
rect 28011 22156 28012 22196
rect 28052 22156 28053 22196
rect 28011 22147 28053 22156
rect 22251 21692 22293 21701
rect 22251 21652 22252 21692
rect 22292 21652 22293 21692
rect 22251 21643 22293 21652
rect 22155 19508 22197 19517
rect 22155 19468 22156 19508
rect 22196 19468 22197 19508
rect 22155 19459 22197 19468
rect 22156 19374 22196 19459
rect 22252 19256 22292 21643
rect 25899 21524 25941 21533
rect 25899 21484 25900 21524
rect 25940 21484 25941 21524
rect 25899 21475 25941 21484
rect 26859 21524 26901 21533
rect 26859 21484 26860 21524
rect 26900 21484 26901 21524
rect 26859 21475 26901 21484
rect 27436 21524 27476 21533
rect 22347 21356 22389 21365
rect 22347 21316 22348 21356
rect 22388 21316 22389 21356
rect 22347 21307 22389 21316
rect 22348 20012 22388 21307
rect 25900 21113 25940 21475
rect 26475 21440 26517 21449
rect 26475 21400 26476 21440
rect 26516 21400 26517 21440
rect 26475 21391 26517 21400
rect 26476 21306 26516 21391
rect 26860 21390 26900 21475
rect 27052 21440 27092 21449
rect 26956 21400 27052 21440
rect 26956 21356 26996 21400
rect 27052 21391 27092 21400
rect 27436 21365 27476 21484
rect 26955 21316 26996 21356
rect 27435 21356 27477 21365
rect 27435 21316 27436 21356
rect 27476 21316 27477 21356
rect 26859 21272 26901 21281
rect 26955 21272 26995 21316
rect 27435 21307 27477 21316
rect 26764 21232 26860 21272
rect 26900 21232 26995 21272
rect 25899 21104 25941 21113
rect 25899 21064 25900 21104
rect 25940 21064 25941 21104
rect 25899 21055 25941 21064
rect 26667 21020 26709 21029
rect 26667 20980 26668 21020
rect 26708 20980 26709 21020
rect 26667 20971 26709 20980
rect 25804 20600 25844 20609
rect 24075 20264 24117 20273
rect 24075 20224 24076 20264
rect 24116 20224 24117 20264
rect 24075 20215 24117 20224
rect 22348 19963 22388 19972
rect 22732 20096 22772 20105
rect 22539 19844 22581 19853
rect 22539 19804 22540 19844
rect 22580 19804 22581 19844
rect 22539 19795 22581 19804
rect 22540 19710 22580 19795
rect 22732 19592 22772 20056
rect 22828 20096 22868 20105
rect 22828 19853 22868 20056
rect 22924 20096 22964 20105
rect 22827 19844 22869 19853
rect 22827 19804 22828 19844
rect 22868 19804 22869 19844
rect 22827 19795 22869 19804
rect 22540 19552 22772 19592
rect 22348 19256 22388 19265
rect 22252 19216 22348 19256
rect 22348 19207 22388 19216
rect 22444 19256 22484 19265
rect 22540 19256 22580 19552
rect 22828 19340 22868 19795
rect 22732 19300 22868 19340
rect 22540 19242 22676 19256
rect 22540 19216 22636 19242
rect 22156 19088 22196 19097
rect 22059 18668 22101 18677
rect 22059 18628 22060 18668
rect 22100 18628 22101 18668
rect 22059 18619 22101 18628
rect 22060 18500 22100 18619
rect 22156 18500 22196 19048
rect 22444 18509 22484 19216
rect 22636 19193 22676 19202
rect 22540 19088 22580 19097
rect 22732 19088 22772 19300
rect 22540 18929 22580 19048
rect 22636 19048 22772 19088
rect 22828 19172 22868 19181
rect 22539 18920 22581 18929
rect 22539 18880 22540 18920
rect 22580 18880 22581 18920
rect 22539 18871 22581 18880
rect 22539 18584 22581 18593
rect 22539 18544 22540 18584
rect 22580 18544 22581 18584
rect 22539 18535 22581 18544
rect 22252 18500 22292 18509
rect 22156 18460 22252 18500
rect 22060 18451 22100 18460
rect 22252 18451 22292 18460
rect 22443 18500 22485 18509
rect 22443 18460 22444 18500
rect 22484 18460 22485 18500
rect 22443 18451 22485 18460
rect 22251 18332 22293 18341
rect 22251 18292 22252 18332
rect 22292 18292 22293 18332
rect 22251 18283 22293 18292
rect 22443 18332 22485 18341
rect 22443 18292 22444 18332
rect 22484 18292 22485 18332
rect 22443 18283 22485 18292
rect 22252 17828 22292 18283
rect 22444 18198 22484 18283
rect 22443 17996 22485 18005
rect 22443 17956 22444 17996
rect 22484 17956 22485 17996
rect 22443 17947 22485 17956
rect 22444 17862 22484 17947
rect 22252 17779 22292 17788
rect 22540 17417 22580 18535
rect 22636 17921 22676 19048
rect 22828 18929 22868 19132
rect 22924 19097 22964 20056
rect 23020 20096 23060 20105
rect 23060 20056 23156 20096
rect 23020 20047 23060 20056
rect 22923 19088 22965 19097
rect 22923 19048 22924 19088
rect 22964 19048 22965 19088
rect 22923 19039 22965 19048
rect 22827 18920 22869 18929
rect 22827 18880 22828 18920
rect 22868 18880 22869 18920
rect 22827 18871 22869 18880
rect 22924 18761 22964 19039
rect 22923 18752 22965 18761
rect 22923 18712 22924 18752
rect 22964 18712 22965 18752
rect 22923 18703 22965 18712
rect 23116 18677 23156 20056
rect 23308 19928 23348 19937
rect 23212 19888 23308 19928
rect 23212 19256 23252 19888
rect 23308 19879 23348 19888
rect 23212 19207 23252 19216
rect 24076 19256 24116 20215
rect 25612 20021 25652 20106
rect 25804 20105 25844 20560
rect 25803 20096 25845 20105
rect 26668 20096 26708 20971
rect 25803 20056 25804 20096
rect 25844 20056 25845 20096
rect 25803 20047 25845 20056
rect 26476 20056 26668 20096
rect 25611 20012 25653 20021
rect 25611 19972 25612 20012
rect 25652 19972 25653 20012
rect 25611 19963 25653 19972
rect 26283 20012 26325 20021
rect 26283 19972 26284 20012
rect 26324 19972 26325 20012
rect 26283 19963 26325 19972
rect 26284 19878 26324 19963
rect 26476 19928 26516 20056
rect 26668 20047 26708 20056
rect 26764 20021 26804 21232
rect 26859 21223 26901 21232
rect 26860 21138 26900 21223
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 26956 20768 26996 20777
rect 26956 20273 26996 20728
rect 26955 20264 26997 20273
rect 26955 20224 26956 20264
rect 26996 20224 26997 20264
rect 26955 20215 26997 20224
rect 27243 20264 27285 20273
rect 27243 20224 27244 20264
rect 27284 20224 27285 20264
rect 27243 20215 27285 20224
rect 26860 20096 26900 20105
rect 26763 20012 26805 20021
rect 26763 19972 26764 20012
rect 26804 19972 26805 20012
rect 26763 19963 26805 19972
rect 26476 19879 26516 19888
rect 25420 19844 25460 19853
rect 26668 19844 26708 19853
rect 25460 19804 25652 19844
rect 25420 19795 25460 19804
rect 23115 18668 23157 18677
rect 23115 18628 23116 18668
rect 23156 18628 23157 18668
rect 23115 18619 23157 18628
rect 22732 18584 22772 18593
rect 22732 18005 22772 18544
rect 23019 18584 23061 18593
rect 23019 18544 23020 18584
rect 23060 18544 23061 18584
rect 23019 18535 23061 18544
rect 22827 18500 22869 18509
rect 22827 18460 22828 18500
rect 22868 18460 22869 18500
rect 22827 18451 22869 18460
rect 22731 17996 22773 18005
rect 22731 17956 22732 17996
rect 22772 17956 22773 17996
rect 22731 17947 22773 17956
rect 22635 17912 22677 17921
rect 22635 17872 22636 17912
rect 22676 17872 22677 17912
rect 22635 17863 22677 17872
rect 22828 17753 22868 18451
rect 23020 18450 23060 18535
rect 23116 18534 23156 18619
rect 23596 18500 23636 18509
rect 23404 18332 23444 18341
rect 23019 18164 23061 18173
rect 23019 18124 23020 18164
rect 23060 18124 23061 18164
rect 23019 18115 23061 18124
rect 22635 17744 22677 17753
rect 22635 17704 22636 17744
rect 22676 17704 22677 17744
rect 22635 17695 22677 17704
rect 22827 17744 22869 17753
rect 22827 17704 22828 17744
rect 22868 17704 22869 17744
rect 22827 17695 22869 17704
rect 22924 17744 22964 17753
rect 22636 17610 22676 17695
rect 22731 17660 22773 17669
rect 22731 17620 22732 17660
rect 22772 17620 22773 17660
rect 22731 17611 22773 17620
rect 22732 17526 22772 17611
rect 22828 17610 22868 17695
rect 22539 17408 22581 17417
rect 22539 17368 22540 17408
rect 22580 17368 22581 17408
rect 22539 17359 22581 17368
rect 22731 17408 22773 17417
rect 22731 17368 22732 17408
rect 22772 17368 22773 17408
rect 22731 17359 22773 17368
rect 22732 17072 22772 17359
rect 22924 17300 22964 17704
rect 22828 17260 22964 17300
rect 23020 17300 23060 18115
rect 23211 17744 23253 17753
rect 23211 17704 23212 17744
rect 23252 17704 23253 17744
rect 23211 17695 23253 17704
rect 23115 17660 23157 17669
rect 23115 17620 23116 17660
rect 23156 17620 23157 17660
rect 23115 17611 23157 17620
rect 23116 17526 23156 17611
rect 23020 17260 23156 17300
rect 22828 17156 22868 17260
rect 22828 17107 22868 17116
rect 22732 17023 22772 17032
rect 22923 17072 22965 17081
rect 22923 17032 22924 17072
rect 22964 17032 22965 17072
rect 22923 17023 22965 17032
rect 23116 17072 23156 17260
rect 23212 17156 23252 17695
rect 23404 17300 23444 18292
rect 23596 18089 23636 18460
rect 23787 18500 23829 18509
rect 23787 18460 23788 18500
rect 23828 18460 23829 18500
rect 23787 18451 23829 18460
rect 23979 18500 24021 18509
rect 23979 18460 23980 18500
rect 24020 18460 24021 18500
rect 23979 18451 24021 18460
rect 23788 18416 23828 18451
rect 23788 18365 23828 18376
rect 23980 18366 24020 18451
rect 23595 18080 23637 18089
rect 23595 18040 23596 18080
rect 23636 18040 23637 18080
rect 23595 18031 23637 18040
rect 23212 17107 23252 17116
rect 23308 17260 23444 17300
rect 23500 17744 23540 17753
rect 24076 17744 24116 19216
rect 25228 19088 25268 19097
rect 25228 18677 25268 19048
rect 25227 18668 25269 18677
rect 25227 18628 25228 18668
rect 25268 18628 25364 18668
rect 25227 18619 25269 18628
rect 25324 18584 25364 18628
rect 25612 18593 25652 19804
rect 25900 19424 25940 19433
rect 25900 19340 25940 19384
rect 25900 19300 26228 19340
rect 26188 19256 26228 19300
rect 26476 19256 26516 19265
rect 26188 19216 26476 19256
rect 26476 19207 26516 19216
rect 26668 19181 26708 19804
rect 26092 19172 26132 19181
rect 26092 18752 26132 19132
rect 26667 19172 26709 19181
rect 26667 19132 26668 19172
rect 26708 19132 26709 19172
rect 26667 19123 26709 19132
rect 26092 18703 26132 18712
rect 26571 18752 26613 18761
rect 26571 18712 26572 18752
rect 26612 18712 26613 18752
rect 26571 18703 26613 18712
rect 25324 18535 25364 18544
rect 25420 18584 25460 18593
rect 24364 18500 24404 18511
rect 24364 18425 24404 18460
rect 24363 18416 24405 18425
rect 24363 18376 24364 18416
rect 24404 18376 24405 18416
rect 24363 18367 24405 18376
rect 24172 18332 24212 18341
rect 24172 18173 24212 18292
rect 24556 18332 24596 18341
rect 24171 18164 24213 18173
rect 24171 18124 24172 18164
rect 24212 18124 24213 18164
rect 24171 18115 24213 18124
rect 24172 17921 24212 18115
rect 24556 18089 24596 18292
rect 25420 18089 25460 18544
rect 25611 18584 25653 18593
rect 25611 18544 25612 18584
rect 25652 18544 25653 18584
rect 25611 18535 25653 18544
rect 25900 18584 25940 18593
rect 25612 18416 25652 18425
rect 25900 18416 25940 18544
rect 25996 18584 26036 18593
rect 26188 18584 26228 18593
rect 26380 18584 26420 18593
rect 26036 18544 26132 18584
rect 25996 18535 26036 18544
rect 25652 18376 25940 18416
rect 25612 18367 25652 18376
rect 24555 18080 24597 18089
rect 24555 18040 24556 18080
rect 24596 18040 24597 18080
rect 24555 18031 24597 18040
rect 25419 18080 25461 18089
rect 25419 18040 25420 18080
rect 25460 18040 25461 18080
rect 25419 18031 25461 18040
rect 24171 17912 24213 17921
rect 24171 17872 24172 17912
rect 24212 17872 24213 17912
rect 24171 17863 24213 17872
rect 24364 17744 24404 17753
rect 24076 17704 24364 17744
rect 23500 17300 23540 17704
rect 24364 17695 24404 17704
rect 23500 17260 23732 17300
rect 23116 17023 23156 17032
rect 23308 17072 23348 17260
rect 23308 17023 23348 17032
rect 22924 16938 22964 17023
rect 23692 16904 23732 17260
rect 24556 17081 24596 18031
rect 26092 17996 26132 18544
rect 26228 18544 26380 18584
rect 26188 18535 26228 18544
rect 26380 18535 26420 18544
rect 26476 18584 26516 18593
rect 26476 18173 26516 18544
rect 26572 18584 26612 18703
rect 26572 18535 26612 18544
rect 26667 18584 26709 18593
rect 26667 18544 26668 18584
rect 26708 18544 26709 18584
rect 26667 18535 26709 18544
rect 26668 18450 26708 18535
rect 26764 18248 26804 19963
rect 26860 19937 26900 20056
rect 26955 20096 26997 20105
rect 26955 20056 26956 20096
rect 26996 20056 26997 20096
rect 27244 20096 27284 20215
rect 27532 20096 27572 22147
rect 27915 22112 27957 22121
rect 27915 22072 27916 22112
rect 27956 22072 27957 22112
rect 27915 22063 27957 22072
rect 28203 22112 28245 22121
rect 28203 22072 28204 22112
rect 28244 22072 28245 22112
rect 28203 22063 28245 22072
rect 27627 21776 27669 21785
rect 27627 21736 27628 21776
rect 27668 21736 27669 21776
rect 27627 21727 27669 21736
rect 27628 21440 27668 21727
rect 27820 21608 27860 21617
rect 27628 21391 27668 21400
rect 27724 21568 27820 21608
rect 27627 20936 27669 20945
rect 27627 20896 27628 20936
rect 27668 20896 27669 20936
rect 27627 20887 27669 20896
rect 27628 20273 27668 20887
rect 27627 20264 27669 20273
rect 27627 20224 27628 20264
rect 27668 20224 27669 20264
rect 27627 20215 27669 20224
rect 27724 20105 27764 21568
rect 27820 21559 27860 21568
rect 27916 21608 27956 22063
rect 28204 21978 28244 22063
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 28779 21944 28821 21953
rect 28779 21904 28780 21944
rect 28820 21904 28821 21944
rect 28779 21895 28821 21904
rect 28011 21776 28053 21785
rect 28011 21736 28012 21776
rect 28052 21736 28053 21776
rect 28011 21727 28053 21736
rect 27916 21559 27956 21568
rect 28012 21608 28052 21727
rect 28395 21692 28437 21701
rect 28395 21652 28396 21692
rect 28436 21652 28437 21692
rect 28395 21643 28437 21652
rect 28012 21559 28052 21568
rect 28108 21608 28148 21617
rect 28300 21608 28340 21617
rect 28148 21568 28300 21608
rect 28108 21559 28148 21568
rect 28300 21559 28340 21568
rect 27819 21440 27861 21449
rect 27819 21400 27820 21440
rect 27860 21400 27861 21440
rect 27819 21391 27861 21400
rect 27820 20768 27860 21391
rect 28300 21356 28340 21365
rect 28011 20852 28053 20861
rect 28011 20812 28012 20852
rect 28052 20812 28053 20852
rect 28011 20803 28053 20812
rect 27820 20719 27860 20728
rect 27915 20684 27957 20693
rect 27915 20644 27916 20684
rect 27956 20644 27957 20684
rect 27915 20635 27957 20644
rect 27723 20096 27765 20105
rect 27244 20056 27476 20096
rect 27532 20056 27668 20096
rect 26955 20047 26997 20056
rect 26956 19962 26996 20047
rect 27148 20012 27188 20021
rect 27436 20012 27476 20056
rect 27436 19972 27572 20012
rect 26859 19928 26901 19937
rect 26859 19888 26860 19928
rect 26900 19888 26901 19928
rect 26859 19879 26901 19888
rect 27148 19844 27188 19972
rect 27339 19928 27381 19937
rect 27339 19888 27340 19928
rect 27380 19888 27381 19928
rect 27339 19879 27381 19888
rect 26956 19804 27188 19844
rect 26956 19760 26996 19804
rect 27340 19794 27380 19879
rect 26860 19720 26996 19760
rect 26860 18425 26900 19720
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 27373 19256 27413 19265
rect 27373 19088 27413 19216
rect 27532 19088 27572 19972
rect 27628 19349 27668 20056
rect 27723 20056 27724 20096
rect 27764 20056 27765 20096
rect 27723 20047 27765 20056
rect 27916 20096 27956 20635
rect 27916 19517 27956 20056
rect 27915 19508 27957 19517
rect 27915 19468 27916 19508
rect 27956 19468 27957 19508
rect 27915 19459 27957 19468
rect 27627 19340 27669 19349
rect 27627 19300 27628 19340
rect 27668 19300 27669 19340
rect 27627 19291 27669 19300
rect 27373 19048 27860 19088
rect 27051 18752 27093 18761
rect 27051 18712 27052 18752
rect 27092 18712 27093 18752
rect 27051 18703 27093 18712
rect 26955 18584 26997 18593
rect 26955 18544 26956 18584
rect 26996 18544 26997 18584
rect 26955 18535 26997 18544
rect 26859 18416 26901 18425
rect 26859 18376 26860 18416
rect 26900 18376 26901 18416
rect 26859 18367 26901 18376
rect 26764 18208 26900 18248
rect 26475 18164 26517 18173
rect 26475 18124 26476 18164
rect 26516 18124 26517 18164
rect 26475 18115 26517 18124
rect 26476 17996 26516 18005
rect 26092 17956 26476 17996
rect 26379 17828 26421 17837
rect 26379 17788 26380 17828
rect 26420 17788 26421 17828
rect 26379 17779 26421 17788
rect 26380 17744 26420 17779
rect 26380 17693 26420 17704
rect 25515 17660 25557 17669
rect 25515 17620 25516 17660
rect 25556 17620 25557 17660
rect 25515 17611 25557 17620
rect 25516 17576 25556 17611
rect 25516 17417 25556 17536
rect 25515 17408 25557 17417
rect 25515 17368 25516 17408
rect 25556 17368 25557 17408
rect 25515 17359 25557 17368
rect 26476 17081 26516 17956
rect 26764 17912 26804 17921
rect 26572 17872 26764 17912
rect 26572 17744 26612 17872
rect 26764 17863 26804 17872
rect 26572 17695 26612 17704
rect 26763 17576 26805 17585
rect 26763 17536 26764 17576
rect 26804 17536 26805 17576
rect 26763 17527 26805 17536
rect 24555 17072 24597 17081
rect 24555 17032 24556 17072
rect 24596 17032 24597 17072
rect 24555 17023 24597 17032
rect 26475 17072 26517 17081
rect 26475 17032 26476 17072
rect 26516 17032 26517 17072
rect 26475 17023 26517 17032
rect 26764 17072 26804 17527
rect 26860 17417 26900 18208
rect 26956 17744 26996 18535
rect 27052 18425 27092 18703
rect 27051 18416 27093 18425
rect 27051 18376 27052 18416
rect 27092 18376 27093 18416
rect 27051 18367 27093 18376
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 27435 17996 27477 18005
rect 27435 17956 27436 17996
rect 27476 17956 27477 17996
rect 27435 17947 27477 17956
rect 27052 17744 27092 17753
rect 26956 17704 27052 17744
rect 27052 17695 27092 17704
rect 27148 17744 27188 17753
rect 26859 17408 26901 17417
rect 26859 17368 26860 17408
rect 26900 17368 26901 17408
rect 26859 17359 26901 17368
rect 27148 17324 27188 17704
rect 27436 17744 27476 17947
rect 27724 17912 27764 17921
rect 27436 17695 27476 17704
rect 27628 17872 27724 17912
rect 27148 17300 27380 17324
rect 27148 17284 27476 17300
rect 27340 17260 27476 17284
rect 26860 17240 26900 17249
rect 26900 17200 27284 17240
rect 26860 17191 26900 17200
rect 27244 17156 27284 17200
rect 27244 17107 27284 17116
rect 26764 17023 26804 17032
rect 26859 17072 26901 17081
rect 26956 17072 26996 17081
rect 26859 17032 26860 17072
rect 26900 17032 26956 17072
rect 26859 17023 26901 17032
rect 26956 17023 26996 17032
rect 27051 17072 27093 17081
rect 27051 17032 27052 17072
rect 27092 17032 27093 17072
rect 27051 17023 27093 17032
rect 27052 16938 27092 17023
rect 23692 16855 23732 16864
rect 27436 16829 27476 17260
rect 27628 17072 27668 17872
rect 27724 17863 27764 17872
rect 27723 17744 27765 17753
rect 27723 17704 27724 17744
rect 27764 17704 27765 17744
rect 27723 17695 27765 17704
rect 27628 17023 27668 17032
rect 27435 16820 27477 16829
rect 27435 16780 27436 16820
rect 27476 16780 27477 16820
rect 27435 16771 27477 16780
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 27724 16400 27764 17695
rect 27820 17300 27860 19048
rect 28012 18257 28052 20803
rect 28204 20768 28244 20777
rect 28300 20768 28340 21316
rect 28244 20728 28340 20768
rect 28204 20719 28244 20728
rect 28396 20693 28436 21643
rect 28492 21608 28532 21617
rect 28492 20777 28532 21568
rect 28588 21608 28628 21617
rect 28780 21608 28820 21895
rect 28628 21568 28820 21608
rect 28876 21608 28916 21617
rect 28588 21559 28628 21568
rect 28876 21029 28916 21568
rect 29067 21608 29109 21617
rect 29067 21568 29068 21608
rect 29108 21568 29204 21608
rect 29067 21559 29109 21568
rect 29068 21474 29108 21559
rect 28972 21356 29012 21365
rect 28875 21020 28917 21029
rect 28875 20980 28876 21020
rect 28916 20980 28917 21020
rect 28875 20971 28917 20980
rect 28683 20852 28725 20861
rect 28683 20812 28684 20852
rect 28724 20812 28725 20852
rect 28683 20803 28725 20812
rect 28491 20768 28533 20777
rect 28491 20728 28492 20768
rect 28532 20728 28533 20768
rect 28491 20719 28533 20728
rect 28684 20768 28724 20803
rect 28684 20717 28724 20728
rect 28875 20768 28917 20777
rect 28875 20728 28876 20768
rect 28916 20728 28917 20768
rect 28875 20719 28917 20728
rect 28972 20768 29012 21316
rect 29067 21020 29109 21029
rect 29067 20980 29068 21020
rect 29108 20980 29109 21020
rect 29067 20971 29109 20980
rect 28972 20719 29012 20728
rect 28395 20684 28437 20693
rect 28395 20644 28396 20684
rect 28436 20644 28437 20684
rect 28395 20635 28437 20644
rect 28779 20684 28821 20693
rect 28779 20644 28780 20684
rect 28820 20644 28821 20684
rect 28779 20635 28821 20644
rect 28780 20550 28820 20635
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 28203 20180 28245 20189
rect 28203 20140 28204 20180
rect 28244 20140 28245 20180
rect 28203 20131 28245 20140
rect 28204 20096 28244 20131
rect 28204 20045 28244 20056
rect 28299 20096 28341 20105
rect 28780 20096 28820 20105
rect 28299 20056 28300 20096
rect 28340 20056 28341 20096
rect 28299 20047 28341 20056
rect 28588 20056 28780 20096
rect 28300 19962 28340 20047
rect 28588 19928 28628 20056
rect 28780 20047 28820 20056
rect 28876 20096 28916 20719
rect 29068 20189 29108 20971
rect 29067 20180 29109 20189
rect 29067 20140 29068 20180
rect 29108 20140 29109 20180
rect 29067 20131 29109 20140
rect 28876 20047 28916 20056
rect 28983 20109 29023 20118
rect 28983 20012 29023 20069
rect 29067 20012 29109 20021
rect 28983 19972 29068 20012
rect 29108 19972 29109 20012
rect 29067 19963 29109 19972
rect 28588 19879 28628 19888
rect 28492 19088 28532 19097
rect 28532 19048 28820 19088
rect 28492 19039 28532 19048
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 28780 18752 28820 19048
rect 28684 18712 28820 18752
rect 28684 18593 28724 18712
rect 28972 18593 29012 18678
rect 29068 18677 29108 19963
rect 29164 19937 29204 21568
rect 29260 20945 29300 23080
rect 29452 23071 29492 23080
rect 29451 21944 29493 21953
rect 29451 21904 29452 21944
rect 29492 21904 29493 21944
rect 29451 21895 29493 21904
rect 29452 21776 29492 21895
rect 29452 21727 29492 21736
rect 29548 21617 29588 23827
rect 30700 23792 30740 23801
rect 30604 22868 30644 22877
rect 30604 22448 30644 22828
rect 30316 22408 30644 22448
rect 30316 22289 30356 22408
rect 29643 22280 29685 22289
rect 29643 22240 29644 22280
rect 29684 22240 29685 22280
rect 29643 22231 29685 22240
rect 30315 22280 30357 22289
rect 30315 22240 30316 22280
rect 30356 22240 30357 22280
rect 30315 22231 30357 22240
rect 30412 22280 30452 22289
rect 29356 21608 29396 21617
rect 29356 21113 29396 21568
rect 29547 21608 29589 21617
rect 29547 21568 29548 21608
rect 29588 21568 29589 21608
rect 29547 21559 29589 21568
rect 29644 21608 29684 22231
rect 30316 22146 30356 22231
rect 30412 22121 30452 22240
rect 30508 22280 30548 22289
rect 30411 22112 30453 22121
rect 30411 22072 30412 22112
rect 30452 22072 30453 22112
rect 30411 22063 30453 22072
rect 30508 22112 30548 22240
rect 30604 22280 30644 22289
rect 30700 22280 30740 23752
rect 30892 23792 30932 23801
rect 30796 23624 30836 23633
rect 30796 23213 30836 23584
rect 30795 23204 30837 23213
rect 30795 23164 30796 23204
rect 30836 23164 30837 23204
rect 30795 23155 30837 23164
rect 30795 22700 30837 22709
rect 30795 22660 30796 22700
rect 30836 22660 30837 22700
rect 30795 22651 30837 22660
rect 30644 22240 30740 22280
rect 30604 22231 30644 22240
rect 30796 22112 30836 22651
rect 30892 22457 30932 23752
rect 30988 23792 31028 23801
rect 30988 23297 31028 23752
rect 30987 23288 31029 23297
rect 30987 23248 30988 23288
rect 31028 23248 31029 23288
rect 30987 23239 31029 23248
rect 30987 22616 31029 22625
rect 30987 22576 30988 22616
rect 31028 22576 31029 22616
rect 30987 22567 31029 22576
rect 30891 22448 30933 22457
rect 30891 22408 30892 22448
rect 30932 22408 30933 22448
rect 30891 22399 30933 22408
rect 30508 22072 30836 22112
rect 30892 22280 30932 22289
rect 30988 22280 31028 22567
rect 30932 22240 31028 22280
rect 30508 21785 30548 22072
rect 30507 21776 30549 21785
rect 30507 21736 30508 21776
rect 30548 21736 30549 21776
rect 30507 21727 30549 21736
rect 30892 21701 30932 22240
rect 30891 21692 30933 21701
rect 30891 21652 30892 21692
rect 30932 21652 30933 21692
rect 30891 21643 30933 21652
rect 29644 21559 29684 21568
rect 29548 21474 29588 21559
rect 29836 21440 29876 21449
rect 29355 21104 29397 21113
rect 29355 21064 29356 21104
rect 29396 21064 29397 21104
rect 29355 21055 29397 21064
rect 29259 20936 29301 20945
rect 29259 20896 29260 20936
rect 29300 20896 29301 20936
rect 29259 20887 29301 20896
rect 29644 20768 29684 20777
rect 29836 20768 29876 21400
rect 30507 20936 30549 20945
rect 30507 20896 30508 20936
rect 30548 20896 30549 20936
rect 30507 20887 30549 20896
rect 29684 20728 29876 20768
rect 30508 20768 30548 20887
rect 29644 20719 29684 20728
rect 29259 20684 29301 20693
rect 29259 20644 29260 20684
rect 29300 20644 29301 20684
rect 29259 20635 29301 20644
rect 29260 20550 29300 20635
rect 29163 19928 29205 19937
rect 29740 19928 29780 19937
rect 29163 19888 29164 19928
rect 29204 19888 29205 19928
rect 29163 19879 29205 19888
rect 29644 19888 29740 19928
rect 29644 19256 29684 19888
rect 29740 19879 29780 19888
rect 29644 19207 29684 19216
rect 30508 19256 30548 20728
rect 31084 19265 31124 24499
rect 31948 24380 31988 25264
rect 32044 25304 32084 25313
rect 32044 24548 32084 25264
rect 32140 25304 32180 25313
rect 33195 25304 33237 25313
rect 32180 25264 32852 25304
rect 32140 25255 32180 25264
rect 32236 25136 32276 25145
rect 32236 24632 32276 25096
rect 32523 24716 32565 24725
rect 32523 24676 32524 24716
rect 32564 24676 32565 24716
rect 32523 24667 32565 24676
rect 32428 24632 32468 24641
rect 32236 24592 32428 24632
rect 32428 24583 32468 24592
rect 32524 24582 32564 24667
rect 32620 24632 32660 24641
rect 32044 24508 32372 24548
rect 32236 24380 32276 24389
rect 31948 24340 32236 24380
rect 31755 24296 31797 24305
rect 31755 24256 31756 24296
rect 31796 24256 31797 24296
rect 31755 24247 31797 24256
rect 31468 23885 31508 23970
rect 31467 23876 31509 23885
rect 31467 23836 31468 23876
rect 31508 23836 31509 23876
rect 31467 23827 31509 23836
rect 31467 23708 31509 23717
rect 31467 23668 31468 23708
rect 31508 23668 31509 23708
rect 31467 23659 31509 23668
rect 31275 23288 31317 23297
rect 31275 23248 31276 23288
rect 31316 23248 31317 23288
rect 31275 23239 31317 23248
rect 31276 23154 31316 23239
rect 31371 23204 31413 23213
rect 31371 23164 31372 23204
rect 31412 23164 31413 23204
rect 31371 23155 31413 23164
rect 31180 23120 31220 23129
rect 31180 22448 31220 23080
rect 31372 23120 31412 23155
rect 31372 23069 31412 23080
rect 31468 23120 31508 23659
rect 31660 23624 31700 23633
rect 31660 23213 31700 23584
rect 31659 23204 31701 23213
rect 31659 23164 31660 23204
rect 31700 23164 31701 23204
rect 31659 23155 31701 23164
rect 31468 23071 31508 23080
rect 31467 22448 31509 22457
rect 31180 22408 31412 22448
rect 31180 22280 31220 22289
rect 31180 21869 31220 22240
rect 31275 22280 31317 22289
rect 31275 22240 31276 22280
rect 31316 22240 31317 22280
rect 31275 22231 31317 22240
rect 31276 22146 31316 22231
rect 31179 21860 31221 21869
rect 31179 21820 31180 21860
rect 31220 21820 31221 21860
rect 31179 21811 31221 21820
rect 31372 21281 31412 22408
rect 31467 22408 31468 22448
rect 31508 22408 31509 22448
rect 31467 22399 31509 22408
rect 31564 22448 31604 22457
rect 31604 22408 31700 22448
rect 31564 22399 31604 22408
rect 31468 22280 31508 22399
rect 31468 22240 31604 22280
rect 31564 21692 31604 22240
rect 31564 21643 31604 21652
rect 31467 21608 31509 21617
rect 31467 21568 31468 21608
rect 31508 21568 31509 21608
rect 31467 21559 31509 21568
rect 31660 21608 31700 22408
rect 31756 22121 31796 24247
rect 31851 23960 31893 23969
rect 31851 23920 31852 23960
rect 31892 23920 31893 23960
rect 31851 23911 31893 23920
rect 31852 22709 31892 23911
rect 32044 23792 32084 23801
rect 31947 23288 31989 23297
rect 31947 23248 31948 23288
rect 31988 23248 31989 23288
rect 31947 23239 31989 23248
rect 31851 22700 31893 22709
rect 31851 22660 31852 22700
rect 31892 22660 31893 22700
rect 31851 22651 31893 22660
rect 31852 22280 31892 22289
rect 31948 22280 31988 23239
rect 32044 22625 32084 23752
rect 32140 23717 32180 24340
rect 32236 24331 32276 24340
rect 32332 24305 32372 24508
rect 32331 24296 32373 24305
rect 32331 24256 32332 24296
rect 32372 24256 32373 24296
rect 32331 24247 32373 24256
rect 32620 24044 32660 24592
rect 32715 24632 32757 24641
rect 32715 24592 32716 24632
rect 32756 24592 32757 24632
rect 32715 24583 32757 24592
rect 32716 24498 32756 24583
rect 32236 24004 32660 24044
rect 32139 23708 32181 23717
rect 32139 23668 32140 23708
rect 32180 23668 32181 23708
rect 32139 23659 32181 23668
rect 32236 23540 32276 24004
rect 32812 23969 32852 25264
rect 33195 25264 33196 25304
rect 33236 25264 33237 25304
rect 33195 25255 33237 25264
rect 33388 25304 33428 25313
rect 33196 25170 33236 25255
rect 33292 25136 33332 25145
rect 33292 24641 33332 25096
rect 33291 24632 33333 24641
rect 33291 24592 33292 24632
rect 33332 24592 33333 24632
rect 33291 24583 33333 24592
rect 33388 24389 33428 25264
rect 33484 25304 33524 25927
rect 33579 25892 33621 25901
rect 33579 25852 33580 25892
rect 33620 25852 33621 25892
rect 33579 25843 33621 25852
rect 33484 25255 33524 25264
rect 33580 24557 33620 25843
rect 34252 25304 34292 26179
rect 34347 26144 34389 26153
rect 34347 26104 34348 26144
rect 34388 26104 34389 26144
rect 34347 26095 34389 26104
rect 34636 26144 34676 26153
rect 34348 26010 34388 26095
rect 34636 25985 34676 26104
rect 34731 26144 34773 26153
rect 34731 26104 34732 26144
rect 34772 26104 34773 26144
rect 34731 26095 34773 26104
rect 34635 25976 34677 25985
rect 34635 25936 34636 25976
rect 34676 25936 34677 25976
rect 34635 25927 34677 25936
rect 34732 25556 34772 26095
rect 34732 25507 34772 25516
rect 34252 25255 34292 25264
rect 34348 25304 34388 25313
rect 34348 24716 34388 25264
rect 34444 25304 34484 25313
rect 34444 24800 34484 25264
rect 34540 25304 34580 25313
rect 34732 25304 34772 25313
rect 34580 25264 34732 25304
rect 34540 25255 34580 25264
rect 34732 25255 34772 25264
rect 34635 25136 34677 25145
rect 34635 25096 34636 25136
rect 34676 25096 34677 25136
rect 34635 25087 34677 25096
rect 34444 24760 34580 24800
rect 34348 24676 34484 24716
rect 33579 24548 33621 24557
rect 33579 24508 33580 24548
rect 33620 24508 33621 24548
rect 33579 24499 33621 24508
rect 34347 24548 34389 24557
rect 34347 24508 34348 24548
rect 34388 24508 34389 24548
rect 34347 24499 34389 24508
rect 33195 24380 33237 24389
rect 33195 24340 33196 24380
rect 33236 24340 33237 24380
rect 33195 24331 33237 24340
rect 33387 24380 33429 24389
rect 33387 24340 33388 24380
rect 33428 24340 33429 24380
rect 33387 24331 33429 24340
rect 32716 23960 32756 23969
rect 32524 23920 32716 23960
rect 32331 23792 32373 23801
rect 32331 23752 32332 23792
rect 32372 23752 32373 23792
rect 32331 23743 32373 23752
rect 32332 23658 32372 23743
rect 32428 23717 32468 23802
rect 32427 23708 32469 23717
rect 32427 23668 32428 23708
rect 32468 23668 32469 23708
rect 32427 23659 32469 23668
rect 32236 23500 32468 23540
rect 32331 23372 32373 23381
rect 32331 23332 32332 23372
rect 32372 23332 32373 23372
rect 32331 23323 32373 23332
rect 32332 23120 32372 23323
rect 32428 23204 32468 23500
rect 32428 23129 32468 23164
rect 32043 22616 32085 22625
rect 32043 22576 32044 22616
rect 32084 22576 32085 22616
rect 32043 22567 32085 22576
rect 32332 22448 32372 23080
rect 32427 23120 32469 23129
rect 32427 23080 32428 23120
rect 32468 23080 32469 23120
rect 32427 23071 32469 23080
rect 32524 23120 32564 23920
rect 32716 23911 32756 23920
rect 32811 23960 32853 23969
rect 32811 23920 32812 23960
rect 32852 23920 32853 23960
rect 32811 23911 32853 23920
rect 33100 23708 33140 23717
rect 32715 23288 32757 23297
rect 32715 23248 32716 23288
rect 32756 23248 32757 23288
rect 32715 23239 32757 23248
rect 32812 23288 32852 23297
rect 33100 23288 33140 23668
rect 32852 23248 33140 23288
rect 32812 23239 32852 23248
rect 32619 23204 32661 23213
rect 32619 23164 32620 23204
rect 32660 23164 32661 23204
rect 32619 23155 32661 23164
rect 32524 23071 32564 23080
rect 32428 23040 32468 23071
rect 32332 22408 32373 22448
rect 32333 22364 32373 22408
rect 32332 22324 32373 22364
rect 31892 22240 31988 22280
rect 32043 22280 32085 22289
rect 32043 22240 32044 22280
rect 32084 22240 32085 22280
rect 31755 22112 31797 22121
rect 31755 22072 31756 22112
rect 31796 22072 31797 22112
rect 31755 22063 31797 22072
rect 31660 21559 31700 21568
rect 31371 21272 31413 21281
rect 31371 21232 31372 21272
rect 31412 21232 31413 21272
rect 31371 21223 31413 21232
rect 31179 20936 31221 20945
rect 31179 20896 31180 20936
rect 31220 20896 31221 20936
rect 31179 20887 31221 20896
rect 31180 20777 31220 20887
rect 31179 20768 31221 20777
rect 31179 20728 31180 20768
rect 31220 20728 31221 20768
rect 31179 20719 31221 20728
rect 31180 20096 31220 20719
rect 31180 20047 31220 20056
rect 31468 20021 31508 21559
rect 31659 21020 31701 21029
rect 31659 20980 31660 21020
rect 31700 20980 31701 21020
rect 31659 20971 31701 20980
rect 31660 20886 31700 20971
rect 31852 20861 31892 22240
rect 32043 22231 32085 22240
rect 32140 22280 32180 22289
rect 32044 22146 32084 22231
rect 31948 22112 31988 22121
rect 31948 22028 31988 22072
rect 32043 22028 32085 22037
rect 31948 21988 32044 22028
rect 32084 21988 32085 22028
rect 32043 21979 32085 21988
rect 32043 21860 32085 21869
rect 32043 21820 32044 21860
rect 32084 21820 32085 21860
rect 32043 21811 32085 21820
rect 32044 21608 32084 21811
rect 32140 21692 32180 22240
rect 32332 21785 32372 22324
rect 32524 22196 32564 22205
rect 32524 22037 32564 22156
rect 32523 22028 32565 22037
rect 32523 21988 32524 22028
rect 32564 21988 32565 22028
rect 32523 21979 32565 21988
rect 32331 21776 32373 21785
rect 32331 21736 32332 21776
rect 32372 21736 32373 21776
rect 32331 21727 32373 21736
rect 32140 21643 32180 21652
rect 32044 21559 32084 21568
rect 32236 21608 32276 21617
rect 32620 21608 32660 23155
rect 32716 23120 32756 23239
rect 33196 23213 33236 24331
rect 34348 23801 34388 24499
rect 34444 24305 34484 24676
rect 34443 24296 34485 24305
rect 34443 24256 34444 24296
rect 34484 24256 34485 24296
rect 34443 24247 34485 24256
rect 33484 23792 33524 23801
rect 33387 23708 33429 23717
rect 33387 23668 33388 23708
rect 33428 23668 33429 23708
rect 33387 23659 33429 23668
rect 33195 23204 33237 23213
rect 33195 23164 33196 23204
rect 33236 23164 33237 23204
rect 33195 23155 33237 23164
rect 32716 23071 32756 23080
rect 32811 23120 32853 23129
rect 32908 23120 32948 23129
rect 32811 23080 32812 23120
rect 32852 23080 32908 23120
rect 32811 23071 32853 23080
rect 32908 23071 32948 23080
rect 33003 23120 33045 23129
rect 33003 23080 33004 23120
rect 33044 23080 33045 23120
rect 33003 23071 33045 23080
rect 33196 23120 33236 23155
rect 33292 23129 33332 23214
rect 33004 22986 33044 23071
rect 33196 23070 33236 23080
rect 33291 23120 33333 23129
rect 33291 23080 33292 23120
rect 33332 23080 33333 23120
rect 33291 23071 33333 23080
rect 33388 23120 33428 23659
rect 33388 23071 33428 23080
rect 33484 23060 33524 23752
rect 34347 23792 34389 23801
rect 34347 23752 34348 23792
rect 34388 23752 34389 23792
rect 34347 23743 34389 23752
rect 34348 23658 34388 23743
rect 34444 23465 34484 24247
rect 34540 23969 34580 24760
rect 34539 23960 34581 23969
rect 34539 23920 34540 23960
rect 34580 23920 34581 23960
rect 34539 23911 34581 23920
rect 34540 23549 34580 23911
rect 34539 23540 34581 23549
rect 34539 23500 34540 23540
rect 34580 23500 34581 23540
rect 34539 23491 34581 23500
rect 34443 23456 34485 23465
rect 34443 23416 34444 23456
rect 34484 23416 34485 23456
rect 34443 23407 34485 23416
rect 33484 23020 33620 23060
rect 33580 22952 33620 23020
rect 33580 22903 33620 22912
rect 32715 22700 32757 22709
rect 32715 22660 32716 22700
rect 32756 22660 32757 22700
rect 32715 22651 32757 22660
rect 32276 21568 32660 21608
rect 31851 20852 31893 20861
rect 31851 20812 31852 20852
rect 31892 20812 31893 20852
rect 31851 20803 31893 20812
rect 32044 20852 32084 20861
rect 31852 20600 31892 20609
rect 31892 20560 31988 20600
rect 31852 20551 31892 20560
rect 31755 20180 31797 20189
rect 31755 20140 31756 20180
rect 31796 20140 31797 20180
rect 31755 20131 31797 20140
rect 31467 20012 31509 20021
rect 31467 19972 31468 20012
rect 31508 19972 31509 20012
rect 31467 19963 31509 19972
rect 31660 19844 31700 19853
rect 31564 19804 31660 19844
rect 30508 19207 30548 19216
rect 31083 19256 31125 19265
rect 31083 19216 31084 19256
rect 31124 19216 31125 19256
rect 31083 19207 31125 19216
rect 29260 19172 29300 19181
rect 29260 18752 29300 19132
rect 31564 18920 31604 19804
rect 31660 19795 31700 19804
rect 31660 19097 31700 19182
rect 31659 19088 31701 19097
rect 31659 19048 31660 19088
rect 31700 19048 31701 19088
rect 31659 19039 31701 19048
rect 31564 18880 31700 18920
rect 29356 18752 29396 18761
rect 29260 18712 29356 18752
rect 29356 18703 29396 18712
rect 29067 18668 29109 18677
rect 29067 18628 29068 18668
rect 29108 18628 29109 18668
rect 29067 18619 29109 18628
rect 29931 18668 29973 18677
rect 29931 18628 29932 18668
rect 29972 18628 29973 18668
rect 29931 18619 29973 18628
rect 30603 18668 30645 18677
rect 30603 18628 30604 18668
rect 30644 18628 30645 18668
rect 30603 18619 30645 18628
rect 28683 18584 28725 18593
rect 28683 18544 28684 18584
rect 28724 18544 28725 18584
rect 28683 18535 28725 18544
rect 28780 18584 28820 18593
rect 28684 18450 28724 18535
rect 28011 18248 28053 18257
rect 28011 18208 28012 18248
rect 28052 18208 28053 18248
rect 28011 18199 28053 18208
rect 28780 18173 28820 18544
rect 28971 18584 29013 18593
rect 28971 18544 28972 18584
rect 29012 18544 29013 18584
rect 28971 18535 29013 18544
rect 29164 18584 29204 18593
rect 28972 18416 29012 18425
rect 29164 18416 29204 18544
rect 29012 18376 29204 18416
rect 29260 18584 29300 18593
rect 28972 18367 29012 18376
rect 29260 18341 29300 18544
rect 29452 18584 29492 18593
rect 29644 18584 29684 18593
rect 29492 18544 29644 18584
rect 29452 18535 29492 18544
rect 29644 18535 29684 18544
rect 29740 18584 29780 18593
rect 29259 18332 29301 18341
rect 29259 18292 29260 18332
rect 29300 18292 29301 18332
rect 29259 18283 29301 18292
rect 28779 18164 28821 18173
rect 28779 18124 28780 18164
rect 28820 18124 28821 18164
rect 28779 18115 28821 18124
rect 27915 18080 27957 18089
rect 27915 18040 27916 18080
rect 27956 18040 27957 18080
rect 27915 18031 27957 18040
rect 27916 17753 27956 18031
rect 29740 17921 29780 18544
rect 29836 18584 29876 18593
rect 29836 18425 29876 18544
rect 29932 18584 29972 18619
rect 29932 18533 29972 18544
rect 30220 18584 30260 18593
rect 30220 18425 30260 18544
rect 30508 18584 30548 18593
rect 29835 18416 29877 18425
rect 29835 18376 29836 18416
rect 29876 18376 29877 18416
rect 29835 18367 29877 18376
rect 30219 18416 30261 18425
rect 30219 18376 30220 18416
rect 30260 18376 30261 18416
rect 30219 18367 30261 18376
rect 29739 17912 29781 17921
rect 29739 17872 29740 17912
rect 29780 17872 29781 17912
rect 29739 17863 29781 17872
rect 27915 17744 27957 17753
rect 27915 17704 27916 17744
rect 27956 17704 27957 17744
rect 27915 17695 27957 17704
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 27820 17260 28532 17300
rect 27819 17072 27861 17081
rect 27819 17032 27820 17072
rect 27860 17032 27861 17072
rect 27819 17023 27861 17032
rect 28492 17072 28532 17260
rect 29163 17240 29205 17249
rect 29163 17200 29164 17240
rect 29204 17200 29205 17240
rect 29163 17191 29205 17200
rect 28492 17023 28532 17032
rect 27436 16360 27764 16400
rect 27436 16316 27476 16360
rect 27353 16276 27476 16316
rect 27353 16247 27393 16276
rect 27353 16198 27393 16207
rect 27531 16232 27573 16241
rect 27531 16192 27532 16232
rect 27572 16192 27573 16232
rect 27531 16183 27573 16192
rect 21963 16148 22005 16157
rect 21963 16108 21964 16148
rect 22004 16108 22005 16148
rect 21963 16099 22005 16108
rect 27435 16148 27477 16157
rect 27435 16108 27436 16148
rect 27476 16108 27477 16148
rect 27435 16099 27477 16108
rect 27436 16014 27476 16099
rect 27532 16098 27572 16183
rect 27820 16157 27860 17023
rect 27819 16148 27861 16157
rect 27819 16108 27820 16148
rect 27860 16108 27861 16148
rect 27819 16099 27861 16108
rect 21579 15980 21621 15989
rect 21579 15940 21580 15980
rect 21620 15940 21621 15980
rect 21579 15931 21621 15940
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 9003 15392 9045 15401
rect 9003 15352 9004 15392
rect 9044 15352 9045 15392
rect 9003 15343 9045 15352
rect 7467 15224 7509 15233
rect 7467 15184 7468 15224
rect 7508 15184 7509 15224
rect 7467 15175 7509 15184
rect 7468 14729 7508 15175
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 7467 14720 7509 14729
rect 7467 14680 7468 14720
rect 7508 14680 7509 14720
rect 7467 14671 7509 14680
rect 7468 14216 7508 14671
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 7468 14167 7508 14176
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 6796 13159 6836 13168
rect 6028 12940 6356 12980
rect 5931 12368 5973 12377
rect 5931 12328 5932 12368
rect 5972 12328 5973 12368
rect 5931 12319 5973 12328
rect 5932 12234 5972 12319
rect 6220 11696 6260 12940
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 7467 12368 7509 12377
rect 7467 12328 7468 12368
rect 7508 12328 7509 12368
rect 7467 12319 7509 12328
rect 7468 11789 7508 12319
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 6028 9512 6068 9521
rect 6220 9512 6260 11656
rect 7372 11780 7412 11789
rect 7372 11621 7412 11740
rect 7467 11780 7509 11789
rect 7467 11740 7468 11780
rect 7508 11740 7509 11780
rect 7467 11731 7509 11740
rect 7371 11612 7413 11621
rect 7371 11572 7372 11612
rect 7412 11572 7413 11612
rect 7371 11563 7413 11572
rect 7179 9764 7221 9773
rect 7179 9724 7180 9764
rect 7220 9724 7221 9764
rect 7179 9715 7221 9724
rect 7180 9680 7220 9715
rect 7180 9629 7220 9640
rect 6068 9472 6260 9512
rect 6028 8000 6068 9472
rect 7180 9260 7220 9269
rect 7180 8681 7220 9220
rect 7179 8672 7221 8681
rect 7179 8632 7180 8672
rect 7220 8632 7221 8672
rect 7179 8623 7221 8632
rect 7468 8168 7508 11731
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 29164 9521 29204 17191
rect 29643 16820 29685 16829
rect 29643 16780 29644 16820
rect 29684 16780 29685 16820
rect 29643 16771 29685 16780
rect 29644 16241 29684 16771
rect 29643 16232 29685 16241
rect 29643 16192 29644 16232
rect 29684 16192 29685 16232
rect 29643 16183 29685 16192
rect 29740 15821 29780 17863
rect 29739 15812 29781 15821
rect 29739 15772 29740 15812
rect 29780 15772 29781 15812
rect 29739 15763 29781 15772
rect 29836 15485 29876 18367
rect 30123 18332 30165 18341
rect 30123 18292 30124 18332
rect 30164 18292 30165 18332
rect 30123 18283 30165 18292
rect 29932 17744 29972 17753
rect 29932 17585 29972 17704
rect 30124 17744 30164 18283
rect 30220 18005 30260 18367
rect 30219 17996 30261 18005
rect 30219 17956 30220 17996
rect 30260 17956 30261 17996
rect 30219 17947 30261 17956
rect 30124 17695 30164 17704
rect 30220 17744 30260 17753
rect 30027 17660 30069 17669
rect 30027 17620 30028 17660
rect 30068 17620 30069 17660
rect 30027 17611 30069 17620
rect 29931 17576 29973 17585
rect 29931 17536 29932 17576
rect 29972 17536 29973 17576
rect 29931 17527 29973 17536
rect 30028 17526 30068 17611
rect 30220 17300 30260 17704
rect 30411 17660 30453 17669
rect 30411 17620 30412 17660
rect 30452 17620 30453 17660
rect 30411 17611 30453 17620
rect 30412 17526 30452 17611
rect 30220 17260 30452 17300
rect 30412 16904 30452 17260
rect 30508 17249 30548 18544
rect 30604 18534 30644 18619
rect 31084 18584 31124 18593
rect 30892 18416 30932 18425
rect 31084 18416 31124 18544
rect 31276 18584 31316 18593
rect 31276 18509 31316 18544
rect 31275 18500 31317 18509
rect 31275 18460 31276 18500
rect 31316 18460 31317 18500
rect 31275 18451 31317 18460
rect 30932 18376 31124 18416
rect 30892 18367 30932 18376
rect 31179 18332 31221 18341
rect 31179 18292 31180 18332
rect 31220 18292 31221 18332
rect 31179 18283 31221 18292
rect 31180 18198 31220 18283
rect 31276 17837 31316 18451
rect 31275 17828 31317 17837
rect 31275 17788 31276 17828
rect 31316 17788 31317 17828
rect 31275 17779 31317 17788
rect 31660 17753 31700 18880
rect 31756 18173 31796 20131
rect 31851 19088 31893 19097
rect 31851 19048 31852 19088
rect 31892 19048 31893 19088
rect 31851 19039 31893 19048
rect 31852 18677 31892 19039
rect 31851 18668 31893 18677
rect 31851 18628 31852 18668
rect 31892 18628 31893 18668
rect 31851 18619 31893 18628
rect 31852 18584 31892 18619
rect 31852 18534 31892 18544
rect 31948 18584 31988 20560
rect 32044 20273 32084 20812
rect 32139 20852 32181 20861
rect 32139 20812 32140 20852
rect 32180 20812 32181 20852
rect 32139 20803 32181 20812
rect 32043 20264 32085 20273
rect 32043 20224 32044 20264
rect 32084 20224 32085 20264
rect 32043 20215 32085 20224
rect 31755 18164 31797 18173
rect 31755 18124 31756 18164
rect 31796 18124 31797 18164
rect 31755 18115 31797 18124
rect 30796 17744 30836 17753
rect 30796 17300 30836 17704
rect 31659 17744 31701 17753
rect 31659 17704 31660 17744
rect 31700 17704 31701 17744
rect 31659 17695 31701 17704
rect 31660 17610 31700 17695
rect 31563 17576 31605 17585
rect 31563 17536 31564 17576
rect 31604 17536 31605 17576
rect 31563 17527 31605 17536
rect 30796 17260 30932 17300
rect 30507 17240 30549 17249
rect 30507 17200 30508 17240
rect 30548 17200 30549 17240
rect 30507 17191 30549 17200
rect 30508 17072 30548 17191
rect 30508 17023 30548 17032
rect 30699 17072 30741 17081
rect 30699 17032 30700 17072
rect 30740 17032 30741 17072
rect 30699 17023 30741 17032
rect 30700 16938 30740 17023
rect 30604 16904 30644 16913
rect 30412 16864 30604 16904
rect 30604 16855 30644 16864
rect 30892 16904 30932 17260
rect 30892 16855 30932 16864
rect 31372 16232 31412 16241
rect 31412 16192 31508 16232
rect 31372 16183 31412 16192
rect 30988 16148 31028 16157
rect 30988 15737 31028 16108
rect 30987 15728 31029 15737
rect 30987 15688 30988 15728
rect 31028 15688 31029 15728
rect 30987 15679 31029 15688
rect 29835 15476 29877 15485
rect 29835 15436 29836 15476
rect 29876 15436 29877 15476
rect 29835 15427 29877 15436
rect 31468 15392 31508 16192
rect 31468 15343 31508 15352
rect 30316 14720 30356 14729
rect 31179 14720 31221 14729
rect 30356 14680 30452 14720
rect 30316 14671 30356 14680
rect 29931 14636 29973 14645
rect 29931 14596 29932 14636
rect 29972 14596 29973 14636
rect 29931 14587 29973 14596
rect 29932 14502 29972 14587
rect 30412 13880 30452 14680
rect 31179 14680 31180 14720
rect 31220 14680 31221 14720
rect 31179 14671 31221 14680
rect 31180 14586 31220 14671
rect 31371 14636 31413 14645
rect 31371 14596 31372 14636
rect 31412 14596 31413 14636
rect 31371 14587 31413 14596
rect 31372 13880 31412 14587
rect 31468 14048 31508 14057
rect 31564 14048 31604 17527
rect 31948 17417 31988 18544
rect 32044 20096 32084 20105
rect 31947 17408 31989 17417
rect 31947 17368 31948 17408
rect 31988 17368 31989 17408
rect 31947 17359 31989 17368
rect 31948 17081 31988 17359
rect 31947 17072 31989 17081
rect 31947 17032 31948 17072
rect 31988 17032 31989 17072
rect 31947 17023 31989 17032
rect 32044 15728 32084 20056
rect 32140 19601 32180 20803
rect 32236 20021 32276 21568
rect 32716 21524 32756 22651
rect 32908 22280 32948 22289
rect 33772 22280 33812 22289
rect 32948 22240 33236 22280
rect 32908 22231 32948 22240
rect 32907 22112 32949 22121
rect 32907 22072 32908 22112
rect 32948 22072 32949 22112
rect 32907 22063 32949 22072
rect 32620 21484 32756 21524
rect 32427 21272 32469 21281
rect 32427 21232 32428 21272
rect 32468 21232 32469 21272
rect 32427 21223 32469 21232
rect 32428 21029 32468 21223
rect 32427 21020 32469 21029
rect 32427 20980 32428 21020
rect 32468 20980 32469 21020
rect 32427 20971 32469 20980
rect 32332 20684 32372 20693
rect 32235 20012 32277 20021
rect 32235 19972 32236 20012
rect 32276 19972 32277 20012
rect 32235 19963 32277 19972
rect 32235 19844 32277 19853
rect 32235 19804 32236 19844
rect 32276 19804 32277 19844
rect 32235 19795 32277 19804
rect 32139 19592 32181 19601
rect 32139 19552 32140 19592
rect 32180 19552 32181 19592
rect 32139 19543 32181 19552
rect 32140 19256 32180 19265
rect 32140 18836 32180 19216
rect 32236 19256 32276 19795
rect 32332 19508 32372 20644
rect 32620 20600 32660 21484
rect 32812 21440 32852 21449
rect 32716 21400 32812 21440
rect 32716 20768 32756 21400
rect 32812 21391 32852 21400
rect 32908 21272 32948 22063
rect 33003 21608 33045 21617
rect 33003 21568 33004 21608
rect 33044 21568 33045 21608
rect 33003 21559 33045 21568
rect 32716 20719 32756 20728
rect 32812 21232 32948 21272
rect 32620 20560 32756 20600
rect 32620 20096 32660 20105
rect 32524 20056 32620 20096
rect 32428 19508 32468 19517
rect 32332 19468 32428 19508
rect 32428 19459 32468 19468
rect 32236 19207 32276 19216
rect 32428 19256 32468 19265
rect 32524 19256 32564 20056
rect 32620 20047 32660 20056
rect 32716 20096 32756 20560
rect 32716 20047 32756 20056
rect 32812 20096 32852 21232
rect 33004 20945 33044 21559
rect 33196 21440 33236 22240
rect 33196 21391 33236 21400
rect 33003 20936 33045 20945
rect 33003 20896 33004 20936
rect 33044 20896 33045 20936
rect 33003 20887 33045 20896
rect 32812 20047 32852 20056
rect 32907 20096 32949 20105
rect 32907 20056 32908 20096
rect 32948 20056 32949 20096
rect 32907 20047 32949 20056
rect 32715 19844 32757 19853
rect 32715 19804 32716 19844
rect 32756 19804 32757 19844
rect 32715 19795 32757 19804
rect 32468 19216 32564 19256
rect 32428 19207 32468 19216
rect 32140 18796 32276 18836
rect 32140 18593 32180 18678
rect 32139 18584 32181 18593
rect 32139 18544 32140 18584
rect 32180 18544 32181 18584
rect 32139 18535 32181 18544
rect 32140 18416 32180 18425
rect 32236 18416 32276 18796
rect 32620 18668 32660 18677
rect 32331 18584 32373 18593
rect 32331 18544 32332 18584
rect 32372 18544 32373 18584
rect 32331 18535 32373 18544
rect 32524 18584 32564 18593
rect 32180 18376 32276 18416
rect 32140 18367 32180 18376
rect 32139 18248 32181 18257
rect 32139 18208 32140 18248
rect 32180 18208 32181 18248
rect 32139 18199 32181 18208
rect 31852 15688 32084 15728
rect 32140 15728 32180 18199
rect 32235 17744 32277 17753
rect 32235 17704 32236 17744
rect 32276 17704 32277 17744
rect 32235 17695 32277 17704
rect 32236 16232 32276 17695
rect 32236 16183 32276 16192
rect 32140 15688 32276 15728
rect 31755 15308 31797 15317
rect 31755 15268 31756 15308
rect 31796 15268 31797 15308
rect 31755 15259 31797 15268
rect 31508 14008 31604 14048
rect 31660 14048 31700 14057
rect 31468 13999 31508 14008
rect 31468 13880 31508 13889
rect 31372 13840 31468 13880
rect 30412 13831 30452 13840
rect 31468 13831 31508 13840
rect 31660 13469 31700 14008
rect 31756 14048 31796 15259
rect 31852 14057 31892 15688
rect 31947 15560 31989 15569
rect 31947 15520 31948 15560
rect 31988 15520 31989 15560
rect 31947 15511 31989 15520
rect 32140 15560 32180 15569
rect 31948 15426 31988 15511
rect 32043 15308 32085 15317
rect 32043 15268 32044 15308
rect 32084 15268 32085 15308
rect 32043 15259 32085 15268
rect 32044 15174 32084 15259
rect 32140 14561 32180 15520
rect 32139 14552 32181 14561
rect 32139 14512 32140 14552
rect 32180 14512 32181 14552
rect 32139 14503 32181 14512
rect 32236 14225 32276 15688
rect 32332 15653 32372 18535
rect 32524 18509 32564 18544
rect 32523 18500 32565 18509
rect 32523 18460 32524 18500
rect 32564 18460 32565 18500
rect 32523 18451 32565 18460
rect 32524 17585 32564 18451
rect 32620 18416 32660 18628
rect 32716 18584 32756 19795
rect 32811 19760 32853 19769
rect 32811 19720 32812 19760
rect 32852 19720 32853 19760
rect 32811 19711 32853 19720
rect 32812 19508 32852 19711
rect 32908 19685 32948 20047
rect 32907 19676 32949 19685
rect 32907 19636 32908 19676
rect 32948 19636 32949 19676
rect 32907 19627 32949 19636
rect 33004 19592 33044 20887
rect 33579 20768 33621 20777
rect 33772 20768 33812 22240
rect 34636 21113 34676 25087
rect 34828 23633 34868 26776
rect 35020 26767 35060 26776
rect 34923 26396 34965 26405
rect 34923 26356 34924 26396
rect 34964 26356 34965 26396
rect 34923 26347 34965 26356
rect 34924 26144 34964 26347
rect 35019 26228 35061 26237
rect 35019 26188 35020 26228
rect 35060 26188 35061 26228
rect 35019 26179 35061 26188
rect 34924 26095 34964 26104
rect 35020 26094 35060 26179
rect 35116 25976 35156 26944
rect 34924 25936 35156 25976
rect 35212 26816 35252 26825
rect 35212 25976 35252 26776
rect 35403 26396 35445 26405
rect 35403 26356 35404 26396
rect 35444 26356 35445 26396
rect 35403 26347 35445 26356
rect 35308 25976 35348 25985
rect 35212 25936 35308 25976
rect 34924 25304 34964 25936
rect 35308 25927 35348 25936
rect 35211 25808 35253 25817
rect 35404 25808 35444 26347
rect 35211 25768 35212 25808
rect 35252 25768 35253 25808
rect 35211 25759 35253 25768
rect 35308 25768 35444 25808
rect 35500 26144 35540 26153
rect 35019 25556 35061 25565
rect 35019 25516 35020 25556
rect 35060 25516 35061 25556
rect 35019 25507 35061 25516
rect 34924 25255 34964 25264
rect 35020 25304 35060 25507
rect 35020 25255 35060 25264
rect 35212 24641 35252 25759
rect 35308 25304 35348 25768
rect 35404 25556 35444 25565
rect 35500 25556 35540 26104
rect 35596 26144 35636 26944
rect 38284 26935 38324 26944
rect 36076 26816 36116 26825
rect 35692 26732 35732 26741
rect 35692 26312 35732 26692
rect 35692 26263 35732 26272
rect 35596 26095 35636 26104
rect 35788 26144 35828 26153
rect 35788 25817 35828 26104
rect 36076 25976 36116 26776
rect 36940 26816 36980 26825
rect 36652 26060 36692 26069
rect 36556 26020 36652 26060
rect 36268 25976 36308 25985
rect 36076 25936 36268 25976
rect 36268 25927 36308 25936
rect 35787 25808 35829 25817
rect 35787 25768 35788 25808
rect 35828 25768 35829 25808
rect 35787 25759 35829 25768
rect 35692 25565 35732 25650
rect 35444 25516 35540 25556
rect 35691 25556 35733 25565
rect 35691 25516 35692 25556
rect 35732 25516 35733 25556
rect 35404 25507 35444 25516
rect 35691 25507 35733 25516
rect 35499 25388 35541 25397
rect 35499 25348 35500 25388
rect 35540 25348 35541 25388
rect 35499 25339 35541 25348
rect 35308 25255 35348 25264
rect 35500 25304 35540 25339
rect 35692 25313 35732 25398
rect 35884 25397 35924 25428
rect 35883 25388 35925 25397
rect 35883 25348 35884 25388
rect 35924 25348 35925 25388
rect 35883 25339 35925 25348
rect 35500 25253 35540 25264
rect 35691 25304 35733 25313
rect 35691 25264 35692 25304
rect 35732 25264 35733 25304
rect 35691 25255 35733 25264
rect 35884 25304 35924 25339
rect 35884 25145 35924 25264
rect 35980 25304 36020 25313
rect 35883 25136 35925 25145
rect 35883 25096 35884 25136
rect 35924 25096 35925 25136
rect 35883 25087 35925 25096
rect 35980 24809 36020 25264
rect 36363 25304 36405 25313
rect 36363 25264 36364 25304
rect 36404 25264 36405 25304
rect 36363 25255 36405 25264
rect 35979 24800 36021 24809
rect 35979 24760 35980 24800
rect 36020 24760 36021 24800
rect 35979 24751 36021 24760
rect 35116 24632 35156 24641
rect 35116 24053 35156 24592
rect 35211 24632 35253 24641
rect 35211 24592 35212 24632
rect 35252 24592 35253 24632
rect 35211 24583 35253 24592
rect 35500 24632 35540 24641
rect 35540 24592 35636 24632
rect 35500 24583 35540 24592
rect 35115 24044 35157 24053
rect 35115 24004 35116 24044
rect 35156 24004 35157 24044
rect 35115 23995 35157 24004
rect 34827 23624 34869 23633
rect 34827 23584 34828 23624
rect 34868 23584 34869 23624
rect 34827 23575 34869 23584
rect 35212 23297 35252 24583
rect 35499 24128 35541 24137
rect 35499 24088 35500 24128
rect 35540 24088 35541 24128
rect 35499 24079 35541 24088
rect 35500 24044 35540 24079
rect 35500 23717 35540 24004
rect 35499 23708 35541 23717
rect 35499 23668 35500 23708
rect 35540 23668 35541 23708
rect 35499 23659 35541 23668
rect 35211 23288 35253 23297
rect 35211 23248 35212 23288
rect 35252 23248 35253 23288
rect 35211 23239 35253 23248
rect 35596 23060 35636 24592
rect 35884 24053 35924 24138
rect 35883 24044 35925 24053
rect 35883 24004 35884 24044
rect 35924 24004 35925 24044
rect 35883 23995 35925 24004
rect 35884 23792 35924 23801
rect 35692 23752 35884 23792
rect 35692 23288 35732 23752
rect 35884 23743 35924 23752
rect 35787 23540 35829 23549
rect 35787 23500 35788 23540
rect 35828 23500 35829 23540
rect 35787 23491 35829 23500
rect 35692 23239 35732 23248
rect 35500 23020 35636 23060
rect 35788 23120 35828 23491
rect 35884 23129 35924 23214
rect 35500 22952 35540 23020
rect 35500 22903 35540 22912
rect 35788 22868 35828 23080
rect 35883 23120 35925 23129
rect 35883 23080 35884 23120
rect 35924 23080 35925 23120
rect 35883 23071 35925 23080
rect 35980 23120 36020 24751
rect 36364 24632 36404 25255
rect 36459 25136 36501 25145
rect 36459 25096 36460 25136
rect 36500 25096 36501 25136
rect 36459 25087 36501 25096
rect 36076 23920 36308 23960
rect 36076 23792 36116 23920
rect 36076 23743 36116 23752
rect 36172 23792 36212 23801
rect 36075 23456 36117 23465
rect 36075 23416 36076 23456
rect 36116 23416 36117 23456
rect 36075 23407 36117 23416
rect 36076 23129 36116 23407
rect 36172 23381 36212 23752
rect 36171 23372 36213 23381
rect 36171 23332 36172 23372
rect 36212 23332 36213 23372
rect 36268 23372 36308 23920
rect 36364 23801 36404 24592
rect 36363 23792 36405 23801
rect 36363 23752 36364 23792
rect 36404 23752 36405 23792
rect 36363 23743 36405 23752
rect 36364 23658 36404 23743
rect 36268 23332 36404 23372
rect 36171 23323 36213 23332
rect 36268 23129 36308 23214
rect 36364 23213 36404 23332
rect 36363 23204 36405 23213
rect 36363 23164 36364 23204
rect 36404 23164 36405 23204
rect 36363 23155 36405 23164
rect 35980 23071 36020 23080
rect 36075 23120 36117 23129
rect 36075 23080 36076 23120
rect 36116 23080 36117 23120
rect 36075 23071 36117 23080
rect 36267 23120 36309 23129
rect 36267 23080 36268 23120
rect 36308 23080 36309 23120
rect 36267 23071 36309 23080
rect 35788 22828 36020 22868
rect 34923 22616 34965 22625
rect 34923 22576 34924 22616
rect 34964 22576 34965 22616
rect 34923 22567 34965 22576
rect 34924 22532 34964 22567
rect 34924 22481 34964 22492
rect 35595 22448 35637 22457
rect 35595 22408 35596 22448
rect 35636 22408 35637 22448
rect 35595 22399 35637 22408
rect 35596 22314 35636 22399
rect 35788 22196 35828 22205
rect 34924 22112 34964 22121
rect 34924 21869 34964 22072
rect 34923 21860 34965 21869
rect 34923 21820 34924 21860
rect 34964 21820 34965 21860
rect 34923 21811 34965 21820
rect 35788 21785 35828 22156
rect 35787 21776 35829 21785
rect 35787 21736 35788 21776
rect 35828 21736 35829 21776
rect 35787 21727 35829 21736
rect 35788 21440 35828 21449
rect 34635 21104 34677 21113
rect 34635 21064 34636 21104
rect 34676 21064 34677 21104
rect 34635 21055 34677 21064
rect 33579 20728 33580 20768
rect 33620 20728 33812 20768
rect 33579 20719 33621 20728
rect 33580 20634 33620 20719
rect 33292 20096 33332 20105
rect 33100 20081 33140 20090
rect 33332 20056 33428 20096
rect 33292 20047 33332 20056
rect 33100 19769 33140 20041
rect 33195 19844 33237 19853
rect 33195 19804 33196 19844
rect 33236 19804 33237 19844
rect 33195 19795 33237 19804
rect 33099 19760 33141 19769
rect 33099 19720 33100 19760
rect 33140 19720 33141 19760
rect 33099 19711 33141 19720
rect 33196 19710 33236 19795
rect 33195 19592 33237 19601
rect 33004 19552 33140 19592
rect 32908 19508 32948 19517
rect 32812 19468 32908 19508
rect 32908 19459 32948 19468
rect 33100 19088 33140 19552
rect 33195 19552 33196 19592
rect 33236 19552 33237 19592
rect 33195 19543 33237 19552
rect 33196 19256 33236 19543
rect 33196 19207 33236 19216
rect 33292 19256 33332 19265
rect 33100 19048 33236 19088
rect 32812 18593 32852 18678
rect 32716 18535 32756 18544
rect 32811 18584 32853 18593
rect 33004 18584 33044 18593
rect 32811 18544 32812 18584
rect 32852 18544 32853 18584
rect 32811 18535 32853 18544
rect 32908 18544 33004 18584
rect 32908 18416 32948 18544
rect 33004 18535 33044 18544
rect 32620 18376 32948 18416
rect 32523 17576 32565 17585
rect 32523 17536 32524 17576
rect 32564 17536 32565 17576
rect 32523 17527 32565 17536
rect 32812 17576 32852 17585
rect 32812 17333 32852 17536
rect 33003 17408 33045 17417
rect 33003 17368 33004 17408
rect 33044 17368 33045 17408
rect 33003 17359 33045 17368
rect 32811 17324 32853 17333
rect 32811 17284 32812 17324
rect 32852 17284 32853 17324
rect 32811 17275 32853 17284
rect 32523 16232 32565 16241
rect 32523 16192 32524 16232
rect 32564 16192 32565 16232
rect 32523 16183 32565 16192
rect 32331 15644 32373 15653
rect 32331 15604 32332 15644
rect 32372 15604 32373 15644
rect 32331 15595 32373 15604
rect 32331 14552 32373 14561
rect 32331 14512 32332 14552
rect 32372 14512 32468 14552
rect 32331 14503 32373 14512
rect 32332 14418 32372 14503
rect 32235 14216 32277 14225
rect 32235 14176 32236 14216
rect 32276 14176 32277 14216
rect 32235 14167 32277 14176
rect 32331 14132 32373 14141
rect 32331 14092 32332 14132
rect 32372 14092 32373 14132
rect 32331 14083 32373 14092
rect 31756 13999 31796 14008
rect 31851 14048 31893 14057
rect 31851 14008 31852 14048
rect 31892 14008 31893 14048
rect 31851 13999 31893 14008
rect 31659 13460 31701 13469
rect 31659 13420 31660 13460
rect 31700 13420 31701 13460
rect 31659 13411 31701 13420
rect 31852 13217 31892 13999
rect 32332 13998 32372 14083
rect 32428 14048 32468 14512
rect 32428 13999 32468 14008
rect 32044 13796 32084 13805
rect 32084 13756 32372 13796
rect 32044 13747 32084 13756
rect 31851 13208 31893 13217
rect 31851 13168 31852 13208
rect 31892 13168 31893 13208
rect 31851 13159 31893 13168
rect 32332 13208 32372 13756
rect 32427 13460 32469 13469
rect 32427 13420 32428 13460
rect 32468 13420 32469 13460
rect 32427 13411 32469 13420
rect 32428 13326 32468 13411
rect 32332 13159 32372 13168
rect 32524 13208 32564 16183
rect 32907 15812 32949 15821
rect 32907 15772 32908 15812
rect 32948 15772 32949 15812
rect 32907 15763 32949 15772
rect 32811 15644 32853 15653
rect 32811 15604 32812 15644
rect 32852 15604 32853 15644
rect 32811 15595 32853 15604
rect 32812 15560 32852 15595
rect 32812 15509 32852 15520
rect 32812 15308 32852 15317
rect 32620 15268 32812 15308
rect 32620 13208 32660 15268
rect 32812 15259 32852 15268
rect 32908 14888 32948 15763
rect 33004 15569 33044 17359
rect 33196 16988 33236 19048
rect 33292 18845 33332 19216
rect 33291 18836 33333 18845
rect 33291 18796 33292 18836
rect 33332 18796 33333 18836
rect 33291 18787 33333 18796
rect 33388 18761 33428 20056
rect 33580 19256 33620 19265
rect 33387 18752 33429 18761
rect 33387 18712 33388 18752
rect 33428 18712 33429 18752
rect 33387 18703 33429 18712
rect 33291 18584 33333 18593
rect 33291 18544 33292 18584
rect 33332 18544 33333 18584
rect 33291 18535 33333 18544
rect 33388 18584 33428 18593
rect 33292 17996 33332 18535
rect 33388 18416 33428 18544
rect 33483 18584 33525 18593
rect 33580 18584 33620 19216
rect 33676 18593 33716 20728
rect 34636 20441 34676 21055
rect 35788 20768 35828 21400
rect 35980 21272 36020 22828
rect 36076 21356 36116 23071
rect 36171 22448 36213 22457
rect 36171 22408 36172 22448
rect 36212 22408 36213 22448
rect 36171 22399 36213 22408
rect 36172 22280 36212 22399
rect 36172 22231 36212 22240
rect 36267 21776 36309 21785
rect 36267 21736 36268 21776
rect 36308 21736 36309 21776
rect 36267 21727 36309 21736
rect 36268 21642 36308 21727
rect 36171 21608 36213 21617
rect 36171 21568 36172 21608
rect 36212 21568 36213 21608
rect 36171 21559 36213 21568
rect 36364 21608 36404 23155
rect 36460 22961 36500 25087
rect 36556 23885 36596 26020
rect 36652 26011 36692 26020
rect 36747 25976 36789 25985
rect 36747 25936 36748 25976
rect 36788 25936 36789 25976
rect 36747 25927 36789 25936
rect 36844 25976 36884 25985
rect 36651 24800 36693 24809
rect 36651 24760 36652 24800
rect 36692 24760 36693 24800
rect 36651 24751 36693 24760
rect 36555 23876 36597 23885
rect 36555 23836 36556 23876
rect 36596 23836 36597 23876
rect 36555 23827 36597 23836
rect 36652 23204 36692 24751
rect 36748 24473 36788 25927
rect 36844 25145 36884 25936
rect 36940 25313 36980 26776
rect 38092 26648 38132 26657
rect 38092 26405 38132 26608
rect 38091 26396 38133 26405
rect 38091 26356 38092 26396
rect 38132 26356 38133 26396
rect 38091 26347 38133 26356
rect 38091 26060 38133 26069
rect 38091 26020 38092 26060
rect 38132 26020 38133 26060
rect 38091 26011 38133 26020
rect 37708 25976 37748 25985
rect 37612 25936 37708 25976
rect 37227 25892 37269 25901
rect 37227 25852 37228 25892
rect 37268 25852 37269 25892
rect 37227 25843 37269 25852
rect 36939 25304 36981 25313
rect 36939 25264 36940 25304
rect 36980 25264 36981 25304
rect 36939 25255 36981 25264
rect 37228 25304 37268 25843
rect 37228 25255 37268 25264
rect 37612 25304 37652 25936
rect 37708 25927 37748 25936
rect 38092 25649 38132 26011
rect 38091 25640 38133 25649
rect 38091 25600 38092 25640
rect 38132 25600 38133 25640
rect 38091 25591 38133 25600
rect 37612 25255 37652 25264
rect 38475 25304 38517 25313
rect 38475 25264 38476 25304
rect 38516 25264 38517 25304
rect 38475 25255 38517 25264
rect 38476 25170 38516 25255
rect 36843 25136 36885 25145
rect 36843 25096 36844 25136
rect 36884 25096 36885 25136
rect 36843 25087 36885 25096
rect 37515 24800 37557 24809
rect 37515 24760 37516 24800
rect 37556 24760 37557 24800
rect 37515 24751 37557 24760
rect 37516 24666 37556 24751
rect 37707 24716 37749 24725
rect 37707 24676 37708 24716
rect 37748 24676 37749 24716
rect 37707 24667 37749 24676
rect 36747 24464 36789 24473
rect 36747 24424 36748 24464
rect 36788 24424 36789 24464
rect 36747 24415 36789 24424
rect 36652 23155 36692 23164
rect 36748 23129 36788 24415
rect 37036 23960 37076 23969
rect 36939 23288 36981 23297
rect 36939 23248 36940 23288
rect 36980 23248 36981 23288
rect 36939 23239 36981 23248
rect 36556 23120 36596 23129
rect 36459 22952 36501 22961
rect 36459 22912 36460 22952
rect 36500 22912 36501 22952
rect 36459 22903 36501 22912
rect 36460 22616 36500 22903
rect 36556 22700 36596 23080
rect 36747 23120 36789 23129
rect 36747 23080 36748 23120
rect 36788 23080 36789 23120
rect 36747 23071 36789 23080
rect 36940 22952 36980 23239
rect 37036 23129 37076 23920
rect 37323 23792 37365 23801
rect 37323 23752 37324 23792
rect 37364 23752 37365 23792
rect 37323 23743 37365 23752
rect 37324 23658 37364 23743
rect 37227 23624 37269 23633
rect 37227 23584 37228 23624
rect 37268 23584 37269 23624
rect 37227 23575 37269 23584
rect 37228 23456 37268 23575
rect 37228 23416 37364 23456
rect 37131 23288 37173 23297
rect 37131 23248 37132 23288
rect 37172 23248 37173 23288
rect 37131 23239 37173 23248
rect 37035 23120 37077 23129
rect 37035 23080 37036 23120
rect 37076 23080 37077 23120
rect 37035 23071 37077 23080
rect 37132 23120 37172 23239
rect 37227 23204 37269 23213
rect 37227 23164 37228 23204
rect 37268 23164 37269 23204
rect 37227 23155 37269 23164
rect 37132 23071 37172 23080
rect 36940 22903 36980 22912
rect 36556 22660 36692 22700
rect 36460 22576 36596 22616
rect 36364 21559 36404 21568
rect 36460 21608 36500 21617
rect 36556 21608 36596 22576
rect 36652 22457 36692 22660
rect 36651 22448 36693 22457
rect 36651 22408 36652 22448
rect 36692 22408 36693 22448
rect 36651 22399 36693 22408
rect 36843 22448 36885 22457
rect 36843 22408 36844 22448
rect 36884 22408 36885 22448
rect 36843 22399 36885 22408
rect 36652 21608 36692 21617
rect 36556 21568 36652 21608
rect 36172 21474 36212 21559
rect 36460 21440 36500 21568
rect 36652 21559 36692 21568
rect 36844 21608 36884 22399
rect 37036 22280 37076 23071
rect 37228 23070 37268 23155
rect 37324 23120 37364 23416
rect 37036 22231 37076 22240
rect 36844 21559 36884 21568
rect 36748 21440 36788 21449
rect 36460 21400 36748 21440
rect 36748 21391 36788 21400
rect 36076 21316 36212 21356
rect 35980 21232 36116 21272
rect 35788 20719 35828 20728
rect 35404 20684 35444 20693
rect 34732 20600 34772 20609
rect 34635 20432 34677 20441
rect 34635 20392 34636 20432
rect 34676 20392 34677 20432
rect 34635 20383 34677 20392
rect 34732 20105 34772 20560
rect 35211 20432 35253 20441
rect 35211 20392 35212 20432
rect 35252 20392 35253 20432
rect 35211 20383 35253 20392
rect 34827 20180 34869 20189
rect 34827 20140 34828 20180
rect 34868 20140 34869 20180
rect 34827 20131 34869 20140
rect 35019 20180 35061 20189
rect 35019 20140 35020 20180
rect 35060 20140 35061 20180
rect 35019 20131 35061 20140
rect 34731 20096 34773 20105
rect 34731 20056 34732 20096
rect 34772 20056 34773 20096
rect 34731 20047 34773 20056
rect 34828 20021 34868 20131
rect 34923 20096 34965 20105
rect 34923 20056 34924 20096
rect 34964 20056 34965 20096
rect 34923 20047 34965 20056
rect 35020 20096 35060 20131
rect 34827 20012 34869 20021
rect 34827 19972 34828 20012
rect 34868 19972 34869 20012
rect 34827 19963 34869 19972
rect 34924 19962 34964 20047
rect 35020 19937 35060 20056
rect 35212 20096 35252 20383
rect 35404 20264 35444 20644
rect 35692 20264 35732 20273
rect 35404 20224 35692 20264
rect 35692 20215 35732 20224
rect 35212 20047 35252 20056
rect 35500 20096 35540 20105
rect 35019 19928 35061 19937
rect 35019 19888 35020 19928
rect 35060 19888 35061 19928
rect 35019 19879 35061 19888
rect 35212 19928 35252 19937
rect 35500 19928 35540 20056
rect 35252 19888 35540 19928
rect 35596 20096 35636 20105
rect 35212 19879 35252 19888
rect 35596 19508 35636 20056
rect 35788 20096 35828 20105
rect 35980 20096 36020 20105
rect 35828 20056 35980 20096
rect 35788 20047 35828 20056
rect 35980 20047 36020 20056
rect 36076 20096 36116 21232
rect 36076 20047 36116 20056
rect 36172 20096 36212 21316
rect 37131 20936 37173 20945
rect 37131 20896 37132 20936
rect 37172 20896 37173 20936
rect 37131 20887 37173 20896
rect 36651 20768 36693 20777
rect 36651 20728 36652 20768
rect 36692 20728 36693 20768
rect 36651 20719 36693 20728
rect 36652 20634 36692 20719
rect 36172 20047 36212 20056
rect 36267 20096 36309 20105
rect 36267 20056 36268 20096
rect 36308 20056 36309 20096
rect 36267 20047 36309 20056
rect 35788 19508 35828 19517
rect 35596 19468 35788 19508
rect 33868 19424 33908 19433
rect 33483 18544 33484 18584
rect 33524 18544 33620 18584
rect 33675 18584 33717 18593
rect 33675 18544 33676 18584
rect 33716 18544 33717 18584
rect 33483 18535 33525 18544
rect 33675 18535 33717 18544
rect 33388 18376 33595 18416
rect 33555 18332 33595 18376
rect 33868 18332 33908 19384
rect 35692 19256 35732 19265
rect 35596 19216 35692 19256
rect 35596 18677 35636 19216
rect 35692 19207 35732 19216
rect 35788 19088 35828 19468
rect 36076 19424 36116 19433
rect 35884 19256 35924 19265
rect 36076 19256 36116 19384
rect 35924 19216 36116 19256
rect 36268 19256 36308 20047
rect 36364 19256 36404 19265
rect 36268 19216 36364 19256
rect 35884 19207 35924 19216
rect 36364 19207 36404 19216
rect 36460 19256 36500 19265
rect 35788 19048 35924 19088
rect 34827 18668 34869 18677
rect 34827 18628 34828 18668
rect 34868 18628 34869 18668
rect 34827 18619 34869 18628
rect 35595 18668 35637 18677
rect 35595 18628 35596 18668
rect 35636 18628 35637 18668
rect 35595 18619 35637 18628
rect 35787 18668 35829 18677
rect 35787 18628 35788 18668
rect 35828 18628 35829 18668
rect 35787 18619 35829 18628
rect 34251 18584 34293 18593
rect 34251 18544 34252 18584
rect 34292 18544 34293 18584
rect 34251 18535 34293 18544
rect 34252 18450 34292 18535
rect 33555 18292 33908 18332
rect 33483 18248 33525 18257
rect 33483 18208 33484 18248
rect 33524 18208 33525 18248
rect 33483 18199 33525 18208
rect 33388 17996 33428 18005
rect 33292 17956 33388 17996
rect 33388 17947 33428 17956
rect 33291 17744 33333 17753
rect 33291 17704 33292 17744
rect 33332 17704 33333 17744
rect 33291 17695 33333 17704
rect 33484 17744 33524 18199
rect 33579 18164 33621 18173
rect 33579 18124 33580 18164
rect 33620 18124 33621 18164
rect 33579 18115 33621 18124
rect 33484 17695 33524 17704
rect 33292 17417 33332 17695
rect 33580 17492 33620 18115
rect 34732 17912 34772 17921
rect 34155 17744 34197 17753
rect 34155 17704 34156 17744
rect 34196 17704 34197 17744
rect 34155 17695 34197 17704
rect 34348 17744 34388 17753
rect 34156 17610 34196 17695
rect 34252 17660 34292 17669
rect 33484 17452 33620 17492
rect 33291 17408 33333 17417
rect 33291 17368 33292 17408
rect 33332 17368 33333 17408
rect 33291 17359 33333 17368
rect 33388 16988 33428 16997
rect 33196 16948 33388 16988
rect 33388 16939 33428 16948
rect 33484 16409 33524 17452
rect 34252 17324 34292 17620
rect 34060 17284 34292 17324
rect 33868 17156 33908 17165
rect 33772 17072 33812 17081
rect 33580 16820 33620 16829
rect 33772 16820 33812 17032
rect 33868 16904 33908 17116
rect 33964 17081 34004 17166
rect 33963 17072 34005 17081
rect 33963 17032 33964 17072
rect 34004 17032 34005 17072
rect 33963 17023 34005 17032
rect 34060 17072 34100 17284
rect 34060 17023 34100 17032
rect 34252 17072 34292 17081
rect 34252 16904 34292 17032
rect 34348 16913 34388 17704
rect 34539 17072 34581 17081
rect 34539 17032 34540 17072
rect 34580 17032 34581 17072
rect 34539 17023 34581 17032
rect 34636 17072 34676 17081
rect 34732 17072 34772 17872
rect 34676 17032 34772 17072
rect 34636 17023 34676 17032
rect 33868 16864 34292 16904
rect 34347 16904 34389 16913
rect 34347 16864 34348 16904
rect 34388 16864 34389 16904
rect 34347 16855 34389 16864
rect 33620 16780 33812 16820
rect 33483 16400 33525 16409
rect 33483 16360 33484 16400
rect 33524 16360 33525 16400
rect 33483 16351 33525 16360
rect 33580 16325 33620 16780
rect 33963 16736 34005 16745
rect 33963 16696 33964 16736
rect 34004 16696 34005 16736
rect 33963 16687 34005 16696
rect 33675 16400 33717 16409
rect 33675 16360 33676 16400
rect 33716 16360 33717 16400
rect 33675 16351 33717 16360
rect 33579 16316 33621 16325
rect 33579 16276 33580 16316
rect 33620 16276 33621 16316
rect 33579 16267 33621 16276
rect 33676 16232 33716 16351
rect 33676 16183 33716 16192
rect 33964 16232 34004 16687
rect 34540 16484 34580 17023
rect 34636 16484 34676 16493
rect 34540 16444 34636 16484
rect 34348 16400 34388 16409
rect 34388 16360 34580 16400
rect 34348 16351 34388 16360
rect 33964 16183 34004 16192
rect 34540 16232 34580 16360
rect 34540 16183 34580 16192
rect 34060 16148 34100 16157
rect 33388 16064 33428 16073
rect 34060 16064 34100 16108
rect 33292 16024 33388 16064
rect 33428 16024 34100 16064
rect 33003 15560 33045 15569
rect 33003 15520 33004 15560
rect 33044 15520 33045 15560
rect 33003 15511 33045 15520
rect 33118 15560 33158 15569
rect 33292 15560 33332 16024
rect 33388 16015 33428 16024
rect 34636 15905 34676 16444
rect 34731 16232 34773 16241
rect 34828 16232 34868 18619
rect 35499 18584 35541 18593
rect 35499 18544 35500 18584
rect 35540 18544 35541 18584
rect 35499 18535 35541 18544
rect 35692 18584 35732 18595
rect 35403 18332 35445 18341
rect 35403 18292 35404 18332
rect 35444 18292 35445 18332
rect 35403 18283 35445 18292
rect 35404 18198 35444 18283
rect 35500 17072 35540 18535
rect 35692 18509 35732 18544
rect 35788 18534 35828 18619
rect 35884 18584 35924 19048
rect 36460 18677 36500 19216
rect 36748 19256 36788 19265
rect 37035 19256 37077 19265
rect 36788 19216 36980 19256
rect 36748 19207 36788 19216
rect 36171 18668 36213 18677
rect 36171 18628 36172 18668
rect 36212 18628 36213 18668
rect 36171 18619 36213 18628
rect 36459 18668 36501 18677
rect 36459 18628 36460 18668
rect 36500 18628 36501 18668
rect 36459 18619 36501 18628
rect 36843 18668 36885 18677
rect 36843 18628 36844 18668
rect 36884 18628 36885 18668
rect 36843 18619 36885 18628
rect 35884 18535 35924 18544
rect 35980 18584 36020 18593
rect 36020 18544 36116 18584
rect 35980 18535 36020 18544
rect 35691 18500 35733 18509
rect 35691 18460 35692 18500
rect 35732 18460 35733 18500
rect 35691 18451 35733 18460
rect 36076 18080 36116 18544
rect 36172 18534 36212 18619
rect 36556 18584 36596 18593
rect 36076 18040 36500 18080
rect 36460 17996 36500 18040
rect 36460 17947 36500 17956
rect 36556 17912 36596 18544
rect 36748 17912 36788 17921
rect 36556 17872 36748 17912
rect 36748 17863 36788 17872
rect 36844 17753 36884 18619
rect 36364 17744 36404 17753
rect 36171 17240 36213 17249
rect 36171 17200 36172 17240
rect 36212 17200 36213 17240
rect 36171 17191 36213 17200
rect 35500 17023 35540 17032
rect 34731 16192 34732 16232
rect 34772 16192 34868 16232
rect 34731 16183 34773 16192
rect 34732 16098 34772 16183
rect 34923 16148 34965 16157
rect 34923 16108 34924 16148
rect 34964 16108 34965 16148
rect 34923 16099 34965 16108
rect 35979 16148 36021 16157
rect 35979 16108 35980 16148
rect 36020 16108 36021 16148
rect 35979 16099 36021 16108
rect 33963 15896 34005 15905
rect 33963 15856 33964 15896
rect 34004 15856 34005 15896
rect 33963 15847 34005 15856
rect 34635 15896 34677 15905
rect 34635 15856 34636 15896
rect 34676 15856 34677 15896
rect 34635 15847 34677 15856
rect 33483 15812 33525 15821
rect 33483 15772 33484 15812
rect 33524 15772 33525 15812
rect 33483 15763 33525 15772
rect 33158 15520 33292 15560
rect 33118 15511 33158 15520
rect 33292 15511 33332 15520
rect 33388 15560 33428 15571
rect 33004 15426 33044 15511
rect 33388 15485 33428 15520
rect 33484 15560 33524 15763
rect 33867 15728 33909 15737
rect 33867 15688 33868 15728
rect 33908 15688 33909 15728
rect 33867 15679 33909 15688
rect 33868 15594 33908 15679
rect 33484 15511 33524 15520
rect 33580 15560 33620 15569
rect 33772 15560 33812 15569
rect 33620 15520 33772 15560
rect 33580 15511 33620 15520
rect 33772 15511 33812 15520
rect 33964 15560 34004 15847
rect 34924 15728 34964 16099
rect 34732 15688 34924 15728
rect 34444 15569 34484 15654
rect 34636 15653 34676 15684
rect 34635 15644 34677 15653
rect 34635 15604 34636 15644
rect 34676 15604 34677 15644
rect 34635 15595 34677 15604
rect 33964 15511 34004 15520
rect 34060 15560 34100 15569
rect 33387 15476 33429 15485
rect 33387 15436 33388 15476
rect 33428 15436 33429 15476
rect 33387 15427 33429 15436
rect 34060 15392 34100 15520
rect 34443 15560 34485 15569
rect 34443 15520 34444 15560
rect 34484 15520 34485 15560
rect 34443 15511 34485 15520
rect 34636 15560 34676 15595
rect 34444 15392 34484 15401
rect 34060 15352 34444 15392
rect 34444 15343 34484 15352
rect 33003 15308 33045 15317
rect 33003 15268 33004 15308
rect 33044 15268 33045 15308
rect 33003 15259 33045 15268
rect 32812 14848 32948 14888
rect 32812 14720 32852 14848
rect 33004 14813 33044 15259
rect 33484 14888 33524 14897
rect 33388 14848 33484 14888
rect 33003 14804 33045 14813
rect 32812 14671 32852 14680
rect 32908 14764 33004 14804
rect 33044 14764 33045 14804
rect 32908 14720 32948 14764
rect 33003 14755 33045 14764
rect 32908 14671 32948 14680
rect 33004 14699 33044 14708
rect 32716 14552 32756 14561
rect 32756 14512 32948 14552
rect 32716 14503 32756 14512
rect 32715 14216 32757 14225
rect 32715 14176 32716 14216
rect 32756 14176 32757 14216
rect 32715 14167 32757 14176
rect 32716 14048 32756 14167
rect 32716 13553 32756 14008
rect 32715 13544 32757 13553
rect 32715 13504 32716 13544
rect 32756 13504 32757 13544
rect 32715 13495 32757 13504
rect 32811 13460 32853 13469
rect 32811 13420 32812 13460
rect 32852 13420 32853 13460
rect 32811 13411 32853 13420
rect 32716 13208 32756 13217
rect 32620 13168 32716 13208
rect 32524 13159 32564 13168
rect 32716 13159 32756 13168
rect 32812 13208 32852 13411
rect 32908 13208 32948 14512
rect 33004 14225 33044 14659
rect 33003 14216 33045 14225
rect 33003 14176 33004 14216
rect 33044 14176 33045 14216
rect 33003 14167 33045 14176
rect 33004 14048 33044 14057
rect 33004 13460 33044 14008
rect 33388 14048 33428 14848
rect 33484 14839 33524 14848
rect 34636 14804 34676 15520
rect 34732 15560 34772 15688
rect 34924 15679 34964 15688
rect 34732 15511 34772 15520
rect 35115 15392 35157 15401
rect 35115 15352 35116 15392
rect 35156 15352 35157 15392
rect 35115 15343 35157 15352
rect 34636 14764 34964 14804
rect 34251 14720 34293 14729
rect 34251 14680 34252 14720
rect 34292 14680 34293 14720
rect 34251 14671 34293 14680
rect 33388 13999 33428 14008
rect 34252 14048 34292 14671
rect 34827 14216 34869 14225
rect 34827 14176 34828 14216
rect 34868 14176 34869 14216
rect 34827 14167 34869 14176
rect 34252 13999 34292 14008
rect 33004 13411 33044 13420
rect 33004 13208 33044 13217
rect 32908 13168 33004 13208
rect 32812 13159 32852 13168
rect 33004 13159 33044 13168
rect 34828 13208 34868 14167
rect 34828 13159 34868 13168
rect 34924 13208 34964 14764
rect 34924 13159 34964 13168
rect 35116 13208 35156 15343
rect 35595 14888 35637 14897
rect 35595 14848 35596 14888
rect 35636 14848 35637 14888
rect 35595 14839 35637 14848
rect 35499 14804 35541 14813
rect 35499 14764 35500 14804
rect 35540 14764 35541 14804
rect 35499 14755 35541 14764
rect 35211 14720 35253 14729
rect 35211 14680 35212 14720
rect 35252 14680 35253 14720
rect 35211 14671 35253 14680
rect 35116 13049 35156 13168
rect 35020 13040 35060 13049
rect 34923 12620 34965 12629
rect 34923 12580 34924 12620
rect 34964 12580 34965 12620
rect 34923 12571 34965 12580
rect 33868 12536 33908 12545
rect 33868 11957 33908 12496
rect 34252 12536 34292 12545
rect 33867 11948 33909 11957
rect 33867 11908 33868 11948
rect 33908 11908 33909 11948
rect 33867 11899 33909 11908
rect 34252 11864 34292 12496
rect 34827 11948 34869 11957
rect 34827 11908 34828 11948
rect 34868 11908 34869 11948
rect 34827 11899 34869 11908
rect 34348 11864 34388 11873
rect 34252 11824 34348 11864
rect 34348 11815 34388 11824
rect 34828 11814 34868 11899
rect 34827 11696 34869 11705
rect 34827 11656 34828 11696
rect 34868 11656 34869 11696
rect 34827 11647 34869 11656
rect 34828 11562 34868 11647
rect 34924 11621 34964 12571
rect 35020 12368 35060 13000
rect 35115 13040 35157 13049
rect 35115 13000 35116 13040
rect 35156 13000 35157 13040
rect 35115 12991 35157 13000
rect 35116 12536 35156 12545
rect 35212 12536 35252 14671
rect 35403 14216 35445 14225
rect 35403 14176 35404 14216
rect 35444 14176 35445 14216
rect 35403 14167 35445 14176
rect 35404 14082 35444 14167
rect 35403 13292 35445 13301
rect 35403 13252 35404 13292
rect 35444 13252 35445 13292
rect 35403 13243 35445 13252
rect 35156 12496 35252 12536
rect 35116 12487 35156 12496
rect 35020 12328 35156 12368
rect 35019 12200 35061 12209
rect 35019 12160 35020 12200
rect 35060 12160 35061 12200
rect 35019 12151 35061 12160
rect 35020 11696 35060 12151
rect 35020 11647 35060 11656
rect 35116 11696 35156 12328
rect 35116 11647 35156 11656
rect 35307 11696 35349 11705
rect 35307 11656 35308 11696
rect 35348 11656 35349 11696
rect 35307 11647 35349 11656
rect 35404 11696 35444 13243
rect 34923 11612 34965 11621
rect 34923 11572 34924 11612
rect 34964 11572 34965 11612
rect 34923 11563 34965 11572
rect 35308 11562 35348 11647
rect 35404 11033 35444 11656
rect 35500 11696 35540 14755
rect 35596 14754 35636 14839
rect 35980 14720 36020 16099
rect 36172 16073 36212 17191
rect 36364 17072 36404 17704
rect 36555 17744 36597 17753
rect 36555 17704 36556 17744
rect 36596 17704 36597 17744
rect 36555 17695 36597 17704
rect 36843 17744 36885 17753
rect 36843 17704 36844 17744
rect 36884 17704 36885 17744
rect 36843 17695 36885 17704
rect 36556 17610 36596 17695
rect 36940 17249 36980 19216
rect 37035 19216 37036 19256
rect 37076 19216 37077 19256
rect 37035 19207 37077 19216
rect 37036 19088 37076 19207
rect 36939 17240 36981 17249
rect 36939 17200 36940 17240
rect 36980 17200 36981 17240
rect 36939 17191 36981 17200
rect 36940 17072 36980 17081
rect 37036 17072 37076 19048
rect 37132 17333 37172 20887
rect 37227 20012 37269 20021
rect 37227 19972 37228 20012
rect 37268 19972 37269 20012
rect 37227 19963 37269 19972
rect 37228 19340 37268 19963
rect 37228 19097 37268 19300
rect 37227 19088 37269 19097
rect 37227 19048 37228 19088
rect 37268 19048 37269 19088
rect 37227 19039 37269 19048
rect 37131 17324 37173 17333
rect 37131 17284 37132 17324
rect 37172 17284 37173 17324
rect 37131 17275 37173 17284
rect 37324 17240 37364 23080
rect 37419 20768 37461 20777
rect 37419 20728 37420 20768
rect 37460 20728 37461 20768
rect 37419 20719 37461 20728
rect 37420 18593 37460 20719
rect 37516 20096 37556 20105
rect 37516 19517 37556 20056
rect 37708 20096 37748 24667
rect 38091 23708 38133 23717
rect 38091 23668 38092 23708
rect 38132 23668 38133 23708
rect 38091 23659 38133 23668
rect 37899 23372 37941 23381
rect 37899 23332 37900 23372
rect 37940 23332 37941 23372
rect 37899 23323 37941 23332
rect 37900 23288 37940 23323
rect 37900 23237 37940 23248
rect 37803 23204 37845 23213
rect 37803 23164 37804 23204
rect 37844 23164 37845 23204
rect 37803 23155 37845 23164
rect 37804 23120 37844 23155
rect 37804 23069 37844 23080
rect 37996 23120 38036 23129
rect 37996 22961 38036 23080
rect 38092 23120 38132 23659
rect 38283 23204 38325 23213
rect 38283 23164 38284 23204
rect 38324 23164 38325 23204
rect 38283 23155 38325 23164
rect 38092 23071 38132 23080
rect 37995 22952 38037 22961
rect 37995 22912 37996 22952
rect 38036 22912 38037 22952
rect 37995 22903 38037 22912
rect 38187 22448 38229 22457
rect 38187 22408 38188 22448
rect 38228 22408 38229 22448
rect 38187 22399 38229 22408
rect 38188 22314 38228 22399
rect 38284 21524 38324 23155
rect 38476 23120 38516 23129
rect 38476 22541 38516 23080
rect 38475 22532 38517 22541
rect 38475 22492 38476 22532
rect 38516 22492 38517 22532
rect 38475 22483 38517 22492
rect 38668 21608 38708 36679
rect 54412 36678 54452 36763
rect 54796 36728 54836 36737
rect 54892 36728 54932 37528
rect 55660 37409 55700 37494
rect 55371 37400 55413 37409
rect 55371 37360 55372 37400
rect 55412 37360 55413 37400
rect 55371 37351 55413 37360
rect 55468 37400 55508 37409
rect 54836 36688 54932 36728
rect 54796 36679 54836 36688
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 49131 36056 49173 36065
rect 49131 36016 49132 36056
rect 49172 36016 49173 36056
rect 49131 36007 49173 36016
rect 50475 36056 50517 36065
rect 50475 36016 50476 36056
rect 50516 36016 50517 36056
rect 50475 36007 50517 36016
rect 43947 35972 43989 35981
rect 43947 35932 43948 35972
rect 43988 35932 43989 35972
rect 43947 35923 43989 35932
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 43948 33293 43988 35923
rect 49132 35922 49172 36007
rect 49611 35636 49653 35645
rect 49611 35596 49612 35636
rect 49652 35596 49653 35636
rect 49611 35587 49653 35596
rect 46540 35216 46580 35225
rect 46732 35216 46772 35225
rect 46580 35176 46676 35216
rect 46540 35167 46580 35176
rect 46540 34964 46580 34973
rect 46156 34924 46540 34964
rect 45963 34544 46005 34553
rect 45963 34504 45964 34544
rect 46004 34504 46005 34544
rect 45963 34495 46005 34504
rect 45964 34410 46004 34495
rect 46156 34376 46196 34924
rect 46540 34915 46580 34924
rect 46539 34544 46581 34553
rect 46539 34504 46540 34544
rect 46580 34504 46581 34544
rect 46539 34495 46581 34504
rect 46156 34327 46196 34336
rect 46540 34376 46580 34495
rect 46540 34327 46580 34336
rect 46444 33872 46484 33881
rect 46636 33872 46676 35176
rect 46732 34208 46772 35176
rect 46828 35216 46868 35225
rect 46828 34553 46868 35176
rect 49612 35216 49652 35587
rect 48460 34964 48500 34973
rect 46827 34544 46869 34553
rect 46827 34504 46828 34544
rect 46868 34504 46869 34544
rect 46827 34495 46869 34504
rect 48460 34385 48500 34924
rect 49228 34553 49268 34638
rect 49227 34544 49269 34553
rect 49227 34504 49228 34544
rect 49268 34504 49269 34544
rect 49227 34495 49269 34504
rect 47404 34376 47444 34385
rect 46732 34168 46868 34208
rect 46484 33832 46676 33872
rect 46444 33823 46484 33832
rect 46540 33704 46580 33713
rect 46252 33536 46292 33545
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 43179 33284 43221 33293
rect 43179 33244 43180 33284
rect 43220 33244 43221 33284
rect 43179 33235 43221 33244
rect 43947 33284 43989 33293
rect 43947 33244 43948 33284
rect 43988 33244 43989 33284
rect 43947 33235 43989 33244
rect 42123 33200 42165 33209
rect 42123 33160 42124 33200
rect 42164 33160 42165 33200
rect 42123 33151 42165 33160
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 40588 32024 40628 32033
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 40492 31352 40532 31361
rect 40588 31352 40628 31984
rect 40971 31688 41013 31697
rect 40971 31648 40972 31688
rect 41012 31648 41013 31688
rect 40971 31639 41013 31648
rect 41835 31688 41877 31697
rect 41835 31648 41836 31688
rect 41876 31648 41877 31688
rect 41835 31639 41877 31648
rect 40532 31312 40628 31352
rect 40492 31303 40532 31312
rect 40108 31268 40148 31277
rect 40108 30437 40148 31228
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 40972 30848 41012 31639
rect 40972 30799 41012 30808
rect 41356 31352 41396 31361
rect 40587 30596 40629 30605
rect 40587 30556 40588 30596
rect 40628 30556 40629 30596
rect 40587 30547 40629 30556
rect 41163 30596 41205 30605
rect 41163 30556 41164 30596
rect 41204 30556 41205 30596
rect 41163 30547 41205 30556
rect 40588 30462 40628 30547
rect 41164 30462 41204 30547
rect 40107 30428 40149 30437
rect 40107 30388 40108 30428
rect 40148 30388 40149 30428
rect 40107 30379 40149 30388
rect 40780 30428 40820 30437
rect 40972 30428 41012 30437
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 40587 30176 40629 30185
rect 40587 30136 40588 30176
rect 40628 30136 40629 30176
rect 40587 30127 40629 30136
rect 39531 30092 39573 30101
rect 39531 30052 39532 30092
rect 39572 30052 39573 30092
rect 39531 30043 39573 30052
rect 40588 30092 40628 30127
rect 38956 30008 38996 30017
rect 38860 29968 38956 30008
rect 38860 29168 38900 29968
rect 38956 29959 38996 29968
rect 38860 29119 38900 29128
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 39532 28412 39572 30043
rect 40588 30041 40628 30052
rect 40780 30017 40820 30388
rect 40876 30388 40972 30428
rect 40011 30008 40053 30017
rect 40011 29968 40012 30008
rect 40052 29968 40053 30008
rect 40011 29959 40053 29968
rect 40779 30008 40821 30017
rect 40779 29968 40780 30008
rect 40820 29968 40821 30008
rect 40779 29959 40821 29968
rect 40012 29924 40052 29959
rect 40012 29873 40052 29884
rect 40396 29924 40436 29933
rect 40204 29672 40244 29681
rect 40396 29672 40436 29884
rect 40244 29632 40436 29672
rect 40780 29840 40820 29849
rect 39724 29168 39764 29177
rect 39532 28363 39572 28372
rect 39628 29128 39724 29168
rect 39052 27656 39092 27665
rect 39628 27656 39668 29128
rect 39724 29119 39764 29128
rect 40204 29009 40244 29632
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 40780 29168 40820 29800
rect 40876 29840 40916 30388
rect 40972 30379 41012 30388
rect 41356 30269 41396 31312
rect 41836 30353 41876 31639
rect 41931 31184 41973 31193
rect 41931 31144 41932 31184
rect 41972 31144 41973 31184
rect 41931 31135 41973 31144
rect 41835 30344 41877 30353
rect 41835 30304 41836 30344
rect 41876 30304 41877 30344
rect 41835 30295 41877 30304
rect 40971 30260 41013 30269
rect 40971 30220 40972 30260
rect 41012 30220 41013 30260
rect 40971 30211 41013 30220
rect 41355 30260 41397 30269
rect 41355 30220 41356 30260
rect 41396 30220 41397 30260
rect 41355 30211 41397 30220
rect 40876 29791 40916 29800
rect 40972 29840 41012 30211
rect 41835 30176 41877 30185
rect 41835 30136 41836 30176
rect 41876 30136 41877 30176
rect 41835 30127 41877 30136
rect 41643 30092 41685 30101
rect 41643 30052 41644 30092
rect 41684 30052 41685 30092
rect 41643 30043 41685 30052
rect 41260 29840 41300 29849
rect 40972 29791 41012 29800
rect 41164 29800 41260 29840
rect 41068 29672 41108 29681
rect 40972 29632 41068 29672
rect 40875 29168 40917 29177
rect 40780 29128 40876 29168
rect 40916 29128 40917 29168
rect 40875 29119 40917 29128
rect 40203 29000 40245 29009
rect 40203 28960 40204 29000
rect 40244 28960 40245 29000
rect 40203 28951 40245 28960
rect 40876 28916 40916 29119
rect 40107 28748 40149 28757
rect 40107 28708 40108 28748
rect 40148 28708 40149 28748
rect 40107 28699 40149 28708
rect 40108 28412 40148 28699
rect 40108 28363 40148 28372
rect 40492 28337 40532 28422
rect 39723 28328 39765 28337
rect 40300 28328 40340 28337
rect 39723 28288 39724 28328
rect 39764 28288 39765 28328
rect 39723 28279 39765 28288
rect 40204 28288 40300 28328
rect 39724 28160 39764 28279
rect 39724 28111 39764 28120
rect 39916 28160 39956 28169
rect 39956 28120 40148 28160
rect 39916 28111 39956 28120
rect 38956 27616 39052 27656
rect 39092 27616 39668 27656
rect 38859 26060 38901 26069
rect 38859 26020 38860 26060
rect 38900 26020 38901 26060
rect 38859 26011 38901 26020
rect 38860 25926 38900 26011
rect 38956 25313 38996 27616
rect 39052 27607 39092 27616
rect 39723 27320 39765 27329
rect 39723 27280 39724 27320
rect 39764 27280 39765 27320
rect 39723 27271 39765 27280
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 39147 27068 39189 27077
rect 39147 27028 39148 27068
rect 39188 27028 39189 27068
rect 39147 27019 39189 27028
rect 39724 27068 39764 27271
rect 39724 27019 39764 27028
rect 39915 27068 39957 27077
rect 39915 27028 39916 27068
rect 39956 27028 39957 27068
rect 39915 27019 39957 27028
rect 39148 26900 39188 27019
rect 39340 26984 39380 26995
rect 39340 26909 39380 26944
rect 39148 26851 39188 26860
rect 39339 26900 39381 26909
rect 39339 26860 39340 26900
rect 39380 26860 39381 26900
rect 39339 26851 39381 26860
rect 39531 26900 39573 26909
rect 39531 26860 39532 26900
rect 39572 26860 39573 26900
rect 39531 26851 39573 26860
rect 39532 26766 39572 26851
rect 39916 26816 39956 27019
rect 40012 26825 40052 26910
rect 39051 26732 39093 26741
rect 39051 26692 39052 26732
rect 39092 26692 39093 26732
rect 39051 26683 39093 26692
rect 39052 26321 39092 26683
rect 39724 26648 39764 26657
rect 39916 26648 39956 26776
rect 40011 26816 40053 26825
rect 40011 26776 40012 26816
rect 40052 26776 40053 26816
rect 40011 26767 40053 26776
rect 40108 26816 40148 28120
rect 40204 27581 40244 28288
rect 40300 28279 40340 28288
rect 40491 28328 40533 28337
rect 40491 28288 40492 28328
rect 40532 28288 40533 28328
rect 40491 28279 40533 28288
rect 40588 28328 40628 28337
rect 40876 28328 40916 28876
rect 40628 28288 40916 28328
rect 40972 28328 41012 29632
rect 41068 29623 41108 29632
rect 41068 29000 41108 29009
rect 41164 29000 41204 29800
rect 41260 29791 41300 29800
rect 41451 29840 41493 29849
rect 41451 29800 41452 29840
rect 41492 29800 41493 29840
rect 41451 29791 41493 29800
rect 41644 29840 41684 30043
rect 41644 29791 41684 29800
rect 41836 29840 41876 30127
rect 41836 29791 41876 29800
rect 41932 29840 41972 31135
rect 42027 30932 42069 30941
rect 42027 30892 42028 30932
rect 42068 30892 42069 30932
rect 42027 30883 42069 30892
rect 41932 29791 41972 29800
rect 41355 29756 41397 29765
rect 41355 29716 41356 29756
rect 41396 29716 41397 29756
rect 41355 29707 41397 29716
rect 41356 29622 41396 29707
rect 41452 29706 41492 29791
rect 41740 29672 41780 29681
rect 41548 29632 41740 29672
rect 41356 29177 41396 29262
rect 41355 29168 41397 29177
rect 41355 29128 41356 29168
rect 41396 29128 41397 29168
rect 41355 29119 41397 29128
rect 41452 29168 41492 29177
rect 41108 28960 41204 29000
rect 41068 28951 41108 28960
rect 41355 28916 41397 28925
rect 41355 28876 41356 28916
rect 41396 28876 41397 28916
rect 41355 28867 41397 28876
rect 41259 28832 41301 28841
rect 41259 28792 41260 28832
rect 41300 28792 41301 28832
rect 41259 28783 41301 28792
rect 41067 28580 41109 28589
rect 41067 28540 41068 28580
rect 41108 28540 41109 28580
rect 41067 28531 41109 28540
rect 41068 28446 41108 28531
rect 41068 28328 41108 28337
rect 40972 28288 41068 28328
rect 40588 28279 40628 28288
rect 41068 28279 41108 28288
rect 41260 28328 41300 28783
rect 41260 28279 41300 28288
rect 41356 28328 41396 28867
rect 41452 28748 41492 29128
rect 41548 28925 41588 29632
rect 41740 29623 41780 29632
rect 42028 29336 42068 30883
rect 42124 30605 42164 33151
rect 42988 33116 43028 33125
rect 43180 33116 43220 33235
rect 46252 33140 46292 33496
rect 46540 33140 46580 33664
rect 43028 33076 43220 33116
rect 45867 33116 45909 33125
rect 45867 33076 45868 33116
rect 45908 33076 45909 33116
rect 42988 33067 43028 33076
rect 45867 33067 45909 33076
rect 46156 33100 46292 33140
rect 46348 33100 46580 33140
rect 46636 33704 46676 33713
rect 43948 33032 43988 33041
rect 42219 32948 42261 32957
rect 42219 32908 42220 32948
rect 42260 32908 42261 32948
rect 42219 32899 42261 32908
rect 42795 32948 42837 32957
rect 42795 32908 42796 32948
rect 42836 32908 42837 32948
rect 42795 32899 42837 32908
rect 42220 30857 42260 32899
rect 42796 32814 42836 32899
rect 42412 32192 42452 32201
rect 42315 31604 42357 31613
rect 42315 31564 42316 31604
rect 42356 31564 42357 31604
rect 42315 31555 42357 31564
rect 42219 30848 42261 30857
rect 42219 30808 42220 30848
rect 42260 30808 42261 30848
rect 42219 30799 42261 30808
rect 42123 30596 42165 30605
rect 42123 30556 42124 30596
rect 42164 30556 42165 30596
rect 42123 30547 42165 30556
rect 42316 30008 42356 31555
rect 42412 31184 42452 32152
rect 42508 32192 42548 32201
rect 42508 32033 42548 32152
rect 42604 32192 42644 32201
rect 42507 32024 42549 32033
rect 42507 31984 42508 32024
rect 42548 31984 42549 32024
rect 42507 31975 42549 31984
rect 42604 31856 42644 32152
rect 42508 31816 42644 31856
rect 42700 32192 42740 32201
rect 42508 31697 42548 31816
rect 42700 31772 42740 32152
rect 42604 31732 42740 31772
rect 42892 32192 42932 32201
rect 42507 31688 42549 31697
rect 42507 31648 42508 31688
rect 42548 31648 42549 31688
rect 42507 31639 42549 31648
rect 42507 31184 42549 31193
rect 42412 31144 42508 31184
rect 42548 31144 42549 31184
rect 42507 31135 42549 31144
rect 42508 31050 42548 31135
rect 42507 30848 42549 30857
rect 42507 30808 42508 30848
rect 42548 30808 42549 30848
rect 42507 30799 42549 30808
rect 42411 30596 42453 30605
rect 42411 30556 42412 30596
rect 42452 30556 42453 30596
rect 42411 30547 42453 30556
rect 42124 29924 42164 29933
rect 42164 29884 42260 29924
rect 42124 29875 42164 29884
rect 42123 29756 42165 29765
rect 42123 29716 42124 29756
rect 42164 29716 42165 29756
rect 42123 29707 42165 29716
rect 41740 29296 42068 29336
rect 41643 29168 41685 29177
rect 41643 29128 41644 29168
rect 41684 29128 41685 29168
rect 41643 29119 41685 29128
rect 41740 29168 41780 29296
rect 41740 29119 41780 29128
rect 41547 28916 41589 28925
rect 41547 28876 41548 28916
rect 41588 28876 41589 28916
rect 41547 28867 41589 28876
rect 41452 28708 41588 28748
rect 41451 28580 41493 28589
rect 41451 28540 41452 28580
rect 41492 28540 41493 28580
rect 41451 28531 41493 28540
rect 41356 28279 41396 28288
rect 40396 28160 40436 28169
rect 41355 28160 41397 28169
rect 40436 28120 40820 28160
rect 40396 28111 40436 28120
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 40491 27740 40533 27749
rect 40491 27700 40492 27740
rect 40532 27700 40533 27740
rect 40491 27691 40533 27700
rect 40396 27656 40436 27665
rect 40300 27616 40396 27656
rect 40203 27572 40245 27581
rect 40203 27532 40204 27572
rect 40244 27532 40245 27572
rect 40203 27523 40245 27532
rect 40204 27404 40244 27413
rect 40204 27077 40244 27364
rect 40203 27068 40245 27077
rect 40203 27028 40204 27068
rect 40244 27028 40245 27068
rect 40203 27019 40245 27028
rect 39916 26608 40052 26648
rect 39051 26312 39093 26321
rect 39051 26272 39052 26312
rect 39092 26272 39093 26312
rect 39051 26263 39093 26272
rect 39052 26178 39092 26263
rect 39244 26144 39284 26153
rect 39435 26144 39477 26153
rect 39284 26104 39380 26144
rect 39244 26095 39284 26104
rect 39244 25901 39284 25986
rect 39340 25985 39380 26104
rect 39435 26104 39436 26144
rect 39476 26104 39477 26144
rect 39435 26095 39477 26104
rect 39532 26144 39572 26153
rect 39436 26010 39476 26095
rect 39339 25976 39381 25985
rect 39339 25936 39340 25976
rect 39380 25936 39381 25976
rect 39532 25976 39572 26104
rect 39724 26144 39764 26608
rect 39916 26144 39956 26153
rect 39724 26095 39764 26104
rect 39820 26104 39916 26144
rect 39724 25976 39764 25985
rect 39532 25936 39724 25976
rect 39339 25927 39381 25936
rect 39724 25927 39764 25936
rect 39243 25892 39285 25901
rect 39243 25852 39244 25892
rect 39284 25852 39285 25892
rect 39243 25843 39285 25852
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 39820 25472 39860 26104
rect 39916 26095 39956 26104
rect 40012 26144 40052 26608
rect 40012 26095 40052 26104
rect 40108 25808 40148 26776
rect 40204 26816 40244 26825
rect 40300 26816 40340 27616
rect 40396 27607 40436 27616
rect 40492 27606 40532 27691
rect 40588 27656 40628 27665
rect 40588 27245 40628 27616
rect 40684 27656 40724 27665
rect 40780 27656 40820 28120
rect 41355 28120 41356 28160
rect 41396 28120 41397 28160
rect 41355 28111 41397 28120
rect 40724 27616 40820 27656
rect 41068 27656 41108 27667
rect 40684 27607 40724 27616
rect 41068 27581 41108 27616
rect 41260 27656 41300 27665
rect 41067 27572 41109 27581
rect 41067 27532 41068 27572
rect 41108 27532 41109 27572
rect 41067 27523 41109 27532
rect 41164 27404 41204 27413
rect 41068 27364 41164 27404
rect 41068 27245 41108 27364
rect 41164 27355 41204 27364
rect 40587 27236 40629 27245
rect 40587 27196 40588 27236
rect 40628 27196 40629 27236
rect 40587 27187 40629 27196
rect 41067 27236 41109 27245
rect 41067 27196 41068 27236
rect 41108 27196 41109 27236
rect 41067 27187 41109 27196
rect 40875 27068 40917 27077
rect 40875 27028 40876 27068
rect 40916 27028 40917 27068
rect 40875 27019 40917 27028
rect 40244 26776 40340 26816
rect 40492 26816 40532 26825
rect 40204 26767 40244 26776
rect 40492 26657 40532 26776
rect 40780 26816 40820 26825
rect 40780 26657 40820 26776
rect 40876 26816 40916 27019
rect 40971 26900 41013 26909
rect 40971 26860 40972 26900
rect 41012 26860 41013 26900
rect 40971 26851 41013 26860
rect 40876 26767 40916 26776
rect 40491 26648 40533 26657
rect 40491 26608 40492 26648
rect 40532 26608 40533 26648
rect 40491 26599 40533 26608
rect 40779 26648 40821 26657
rect 40779 26608 40780 26648
rect 40820 26608 40821 26648
rect 40779 26599 40821 26608
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 40779 26480 40821 26489
rect 40779 26440 40780 26480
rect 40820 26440 40821 26480
rect 40779 26431 40821 26440
rect 40587 26312 40629 26321
rect 40587 26272 40588 26312
rect 40628 26272 40629 26312
rect 40587 26263 40629 26272
rect 40780 26312 40820 26431
rect 40780 26263 40820 26272
rect 40588 26178 40628 26263
rect 40299 26144 40341 26153
rect 40299 26104 40300 26144
rect 40340 26104 40341 26144
rect 40299 26095 40341 26104
rect 40203 25976 40245 25985
rect 40203 25936 40204 25976
rect 40244 25936 40245 25976
rect 40203 25927 40245 25936
rect 39532 25432 39860 25472
rect 40012 25768 40148 25808
rect 38955 25304 38997 25313
rect 38955 25264 38956 25304
rect 38996 25264 38997 25304
rect 38955 25255 38997 25264
rect 39532 24800 39572 25432
rect 39820 25304 39860 25313
rect 39628 25136 39668 25145
rect 39820 25136 39860 25264
rect 39916 25304 39956 25315
rect 39916 25229 39956 25264
rect 40012 25304 40052 25768
rect 40204 25640 40244 25927
rect 39915 25220 39957 25229
rect 39915 25180 39916 25220
rect 39956 25180 39957 25220
rect 39915 25171 39957 25180
rect 39668 25096 39860 25136
rect 39628 25087 39668 25096
rect 39820 25052 39860 25096
rect 40012 25052 40052 25264
rect 40108 25600 40244 25640
rect 40108 25304 40148 25600
rect 40300 25556 40340 26095
rect 40395 26060 40437 26069
rect 40395 26020 40396 26060
rect 40436 26020 40437 26060
rect 40395 26011 40437 26020
rect 40875 26060 40917 26069
rect 40875 26020 40876 26060
rect 40916 26020 40917 26060
rect 40875 26011 40917 26020
rect 40972 26060 41012 26851
rect 41068 26153 41108 27187
rect 41164 27068 41204 27077
rect 41260 27068 41300 27616
rect 41204 27028 41300 27068
rect 41164 27019 41204 27028
rect 41356 26816 41396 28111
rect 41452 27824 41492 28531
rect 41548 28328 41588 28708
rect 41644 28580 41684 29119
rect 41739 29000 41781 29009
rect 41739 28960 41740 29000
rect 41780 28960 41781 29000
rect 41739 28951 41781 28960
rect 41740 28673 41780 28951
rect 41739 28664 41781 28673
rect 41739 28624 41740 28664
rect 41780 28624 41781 28664
rect 41739 28615 41781 28624
rect 41644 28531 41684 28540
rect 41548 27833 41588 28288
rect 41740 28328 41780 28615
rect 41836 28589 41876 29296
rect 42027 29168 42069 29177
rect 42027 29128 42028 29168
rect 42068 29128 42069 29168
rect 42027 29119 42069 29128
rect 42124 29168 42164 29707
rect 42028 29034 42068 29119
rect 42124 29093 42164 29128
rect 42123 29084 42165 29093
rect 42123 29044 42124 29084
rect 42164 29044 42165 29084
rect 42123 29035 42165 29044
rect 42124 29004 42164 29035
rect 41835 28580 41877 28589
rect 41835 28540 41836 28580
rect 41876 28540 41877 28580
rect 41835 28531 41877 28540
rect 41931 28496 41973 28505
rect 41931 28456 41932 28496
rect 41972 28456 41973 28496
rect 41931 28447 41973 28456
rect 41740 28279 41780 28288
rect 41932 28328 41972 28447
rect 41932 28279 41972 28288
rect 41452 27775 41492 27784
rect 41547 27824 41589 27833
rect 41547 27784 41548 27824
rect 41588 27784 41589 27824
rect 41547 27775 41589 27784
rect 41644 27572 41684 27581
rect 41644 27413 41684 27532
rect 41452 27404 41492 27413
rect 41452 26909 41492 27364
rect 41643 27404 41685 27413
rect 41643 27364 41644 27404
rect 41684 27364 41685 27404
rect 41643 27355 41685 27364
rect 42220 26984 42260 29884
rect 42316 29849 42356 29968
rect 42315 29840 42357 29849
rect 42315 29800 42316 29840
rect 42356 29800 42357 29840
rect 42315 29791 42357 29800
rect 42315 29168 42357 29177
rect 42315 29128 42316 29168
rect 42356 29128 42357 29168
rect 42315 29119 42357 29128
rect 42316 29034 42356 29119
rect 42316 28916 42356 28925
rect 42316 28505 42356 28876
rect 42412 28757 42452 30547
rect 42508 30176 42548 30799
rect 42604 30596 42644 31732
rect 42892 31688 42932 32152
rect 43084 32192 43124 32201
rect 42700 31648 42932 31688
rect 42988 31940 43028 31949
rect 42700 31604 42740 31648
rect 42700 31555 42740 31564
rect 42988 31445 43028 31900
rect 43084 31613 43124 32152
rect 43276 32192 43316 32201
rect 43660 32192 43700 32201
rect 43948 32192 43988 32992
rect 45676 32864 45716 32873
rect 43316 32152 43604 32192
rect 43276 32143 43316 32152
rect 43564 31688 43604 32152
rect 43700 32152 43988 32192
rect 44524 32192 44564 32201
rect 43660 32143 43700 32152
rect 43564 31648 43988 31688
rect 43083 31604 43125 31613
rect 43083 31564 43084 31604
rect 43124 31564 43125 31604
rect 43083 31555 43125 31564
rect 43948 31604 43988 31648
rect 43948 31555 43988 31564
rect 42987 31436 43029 31445
rect 42892 31396 42988 31436
rect 43028 31396 43029 31436
rect 42892 30680 42932 31396
rect 42987 31387 43029 31396
rect 43084 31352 43124 31361
rect 42988 31268 43028 31279
rect 42988 31193 43028 31228
rect 42987 31184 43029 31193
rect 42987 31144 42988 31184
rect 43028 31144 43029 31184
rect 42987 31135 43029 31144
rect 43084 30848 43124 31312
rect 43372 31352 43412 31361
rect 43660 31352 43700 31361
rect 43372 31025 43412 31312
rect 43468 31312 43660 31352
rect 43371 31016 43413 31025
rect 43371 30976 43372 31016
rect 43412 30976 43413 31016
rect 43371 30967 43413 30976
rect 43468 30848 43508 31312
rect 43660 31303 43700 31312
rect 43755 31352 43797 31361
rect 43948 31352 43988 31361
rect 43755 31312 43756 31352
rect 43796 31312 43797 31352
rect 43755 31303 43797 31312
rect 43852 31312 43948 31352
rect 43756 31218 43796 31303
rect 43084 30808 43316 30848
rect 42988 30680 43028 30689
rect 42796 30669 42836 30678
rect 42892 30640 42988 30680
rect 42988 30631 43028 30640
rect 43084 30680 43124 30689
rect 42796 30596 42836 30629
rect 42604 30556 42836 30596
rect 43084 30521 43124 30640
rect 43276 30680 43316 30808
rect 43372 30808 43508 30848
rect 43372 30764 43412 30808
rect 43372 30715 43412 30724
rect 43276 30605 43316 30640
rect 43468 30680 43508 30689
rect 43275 30596 43317 30605
rect 43275 30556 43276 30596
rect 43316 30556 43317 30596
rect 43275 30547 43317 30556
rect 43083 30512 43125 30521
rect 43083 30472 43084 30512
rect 43124 30472 43125 30512
rect 43083 30463 43125 30472
rect 42604 30428 42644 30439
rect 42604 30353 42644 30388
rect 42795 30428 42837 30437
rect 42795 30388 42796 30428
rect 42836 30388 42837 30428
rect 42795 30379 42837 30388
rect 42603 30344 42645 30353
rect 42603 30304 42604 30344
rect 42644 30304 42645 30344
rect 42603 30295 42645 30304
rect 42796 30294 42836 30379
rect 42508 30136 42644 30176
rect 42508 29000 42548 29009
rect 42411 28748 42453 28757
rect 42411 28708 42412 28748
rect 42452 28708 42453 28748
rect 42411 28699 42453 28708
rect 42315 28496 42357 28505
rect 42315 28456 42316 28496
rect 42356 28456 42357 28496
rect 42315 28447 42357 28456
rect 42316 28328 42356 28337
rect 42508 28328 42548 28960
rect 42356 28288 42548 28328
rect 42316 28279 42356 28288
rect 42028 26944 42260 26984
rect 41451 26900 41493 26909
rect 41451 26860 41452 26900
rect 41492 26860 41493 26900
rect 41451 26851 41493 26860
rect 41260 26776 41356 26816
rect 41067 26144 41109 26153
rect 41067 26104 41068 26144
rect 41108 26104 41109 26144
rect 41067 26095 41109 26104
rect 40972 26011 41012 26020
rect 40396 25926 40436 26011
rect 40588 25892 40628 25901
rect 40779 25892 40821 25901
rect 40628 25852 40724 25892
rect 40588 25843 40628 25852
rect 40396 25556 40436 25565
rect 40300 25516 40396 25556
rect 40300 25304 40340 25313
rect 40108 25255 40148 25264
rect 40204 25264 40300 25304
rect 40107 25136 40149 25145
rect 40107 25096 40108 25136
rect 40148 25096 40149 25136
rect 40107 25087 40149 25096
rect 39820 25012 39956 25052
rect 39532 24760 39668 24800
rect 39532 24632 39572 24641
rect 39051 24548 39093 24557
rect 39051 24508 39052 24548
rect 39092 24508 39093 24548
rect 39051 24499 39093 24508
rect 39052 24414 39092 24499
rect 39244 24389 39284 24474
rect 39532 24473 39572 24592
rect 39531 24464 39573 24473
rect 39531 24424 39532 24464
rect 39572 24424 39573 24464
rect 39531 24415 39573 24424
rect 39243 24380 39285 24389
rect 39243 24340 39244 24380
rect 39284 24340 39285 24380
rect 39243 24331 39285 24340
rect 39628 24305 39668 24760
rect 39820 24632 39860 24643
rect 39820 24557 39860 24592
rect 39916 24632 39956 25012
rect 40011 25012 40052 25052
rect 40011 24968 40051 25012
rect 40011 24928 40052 24968
rect 39819 24548 39861 24557
rect 39819 24508 39820 24548
rect 39860 24508 39861 24548
rect 39819 24499 39861 24508
rect 39627 24296 39669 24305
rect 39532 24256 39628 24296
rect 39668 24256 39669 24296
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 38860 23792 38900 23803
rect 38860 23717 38900 23752
rect 38956 23792 38996 23801
rect 38859 23708 38901 23717
rect 38859 23668 38860 23708
rect 38900 23668 38901 23708
rect 38859 23659 38901 23668
rect 38860 23297 38900 23659
rect 38956 23465 38996 23752
rect 39052 23792 39092 23801
rect 39052 23549 39092 23752
rect 39340 23792 39380 23801
rect 39148 23624 39188 23633
rect 39051 23540 39093 23549
rect 39051 23500 39052 23540
rect 39092 23500 39093 23540
rect 39051 23491 39093 23500
rect 38955 23456 38997 23465
rect 38955 23416 38956 23456
rect 38996 23416 38997 23456
rect 38955 23407 38997 23416
rect 38859 23288 38901 23297
rect 38859 23248 38860 23288
rect 38900 23248 38901 23288
rect 38859 23239 38901 23248
rect 38860 23120 38900 23129
rect 38860 22448 38900 23080
rect 39148 23060 39188 23584
rect 39340 23213 39380 23752
rect 39532 23792 39572 24256
rect 39627 24247 39669 24256
rect 39628 24162 39668 24247
rect 39532 23743 39572 23752
rect 39628 23792 39668 23801
rect 39916 23792 39956 24592
rect 39668 23752 39956 23792
rect 39628 23743 39668 23752
rect 40012 23708 40052 24928
rect 40108 24389 40148 25087
rect 40204 24464 40244 25264
rect 40300 25255 40340 25264
rect 40396 25136 40436 25516
rect 40491 25556 40533 25565
rect 40491 25516 40492 25556
rect 40532 25516 40533 25556
rect 40491 25507 40533 25516
rect 40492 25304 40532 25507
rect 40684 25397 40724 25852
rect 40779 25852 40780 25892
rect 40820 25852 40821 25892
rect 40876 25892 40916 26011
rect 41260 25892 41300 26776
rect 41356 26767 41396 26776
rect 41548 26816 41588 26825
rect 41452 26732 41492 26741
rect 41452 26396 41492 26692
rect 41548 26657 41588 26776
rect 41740 26732 41780 26741
rect 41547 26648 41589 26657
rect 41547 26608 41548 26648
rect 41588 26608 41589 26648
rect 41547 26599 41589 26608
rect 41356 26356 41492 26396
rect 41356 26144 41396 26356
rect 41548 26312 41588 26321
rect 41740 26312 41780 26692
rect 42028 26321 42068 26944
rect 42124 26816 42164 26825
rect 42164 26776 42260 26816
rect 42124 26767 42164 26776
rect 41588 26272 41780 26312
rect 42027 26312 42069 26321
rect 42027 26272 42028 26312
rect 42068 26272 42069 26312
rect 41548 26263 41588 26272
rect 42027 26263 42069 26272
rect 41356 26095 41396 26104
rect 41451 26144 41493 26153
rect 41451 26104 41452 26144
rect 41492 26104 41493 26144
rect 41451 26095 41493 26104
rect 41643 26144 41685 26153
rect 41643 26104 41644 26144
rect 41684 26104 41685 26144
rect 41643 26095 41685 26104
rect 41452 26010 41492 26095
rect 40876 25852 41204 25892
rect 41260 25852 41492 25892
rect 40779 25843 40821 25852
rect 40780 25758 40820 25843
rect 40875 25556 40917 25565
rect 40875 25516 40876 25556
rect 40916 25516 40917 25556
rect 40875 25507 40917 25516
rect 40876 25422 40916 25507
rect 40683 25388 40725 25397
rect 40683 25348 40684 25388
rect 40724 25348 40725 25388
rect 40683 25339 40725 25348
rect 40492 25255 40532 25264
rect 40684 25254 40724 25339
rect 40876 25136 40916 25145
rect 40396 25096 40820 25136
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 40491 24800 40533 24809
rect 40491 24760 40492 24800
rect 40532 24760 40533 24800
rect 40491 24751 40533 24760
rect 40395 24632 40437 24641
rect 40395 24592 40396 24632
rect 40436 24592 40437 24632
rect 40395 24583 40437 24592
rect 40396 24498 40436 24583
rect 40204 24415 40244 24424
rect 40107 24380 40149 24389
rect 40107 24340 40108 24380
rect 40148 24340 40149 24380
rect 40107 24331 40149 24340
rect 40396 24380 40436 24389
rect 39916 23668 40052 23708
rect 39436 23624 39476 23633
rect 39339 23204 39381 23213
rect 39339 23164 39340 23204
rect 39380 23164 39381 23204
rect 39339 23155 39381 23164
rect 38860 22399 38900 22408
rect 38956 23020 39188 23060
rect 39436 23060 39476 23584
rect 39724 23129 39764 23214
rect 39723 23120 39765 23129
rect 39723 23080 39724 23120
rect 39764 23080 39765 23120
rect 39723 23071 39765 23080
rect 39436 23020 39572 23060
rect 38956 22280 38996 23020
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 39051 22532 39093 22541
rect 39051 22492 39052 22532
rect 39092 22492 39093 22532
rect 39051 22483 39093 22492
rect 39052 22398 39092 22483
rect 39052 22280 39092 22289
rect 38956 22240 39052 22280
rect 39052 22231 39092 22240
rect 39243 22280 39285 22289
rect 39243 22240 39244 22280
rect 39284 22240 39285 22280
rect 39243 22231 39285 22240
rect 39340 22280 39380 22289
rect 39532 22280 39572 23020
rect 39380 22240 39572 22280
rect 39340 22231 39380 22240
rect 39244 22146 39284 22231
rect 39052 21608 39092 21617
rect 38668 21568 38804 21608
rect 38188 21484 38324 21524
rect 37804 20600 37844 20609
rect 37804 20105 37844 20560
rect 38188 20441 38228 21484
rect 38571 21356 38613 21365
rect 38571 21316 38572 21356
rect 38612 21316 38613 21356
rect 38571 21307 38613 21316
rect 38284 20768 38324 20777
rect 38187 20432 38229 20441
rect 38187 20392 38188 20432
rect 38228 20392 38229 20432
rect 38187 20383 38229 20392
rect 37708 20047 37748 20056
rect 37803 20096 37845 20105
rect 37900 20096 37940 20105
rect 37803 20056 37804 20096
rect 37844 20056 37900 20096
rect 37803 20047 37845 20056
rect 37900 20047 37940 20056
rect 37995 20096 38037 20105
rect 37995 20056 37996 20096
rect 38036 20056 38037 20096
rect 37995 20047 38037 20056
rect 38188 20096 38228 20383
rect 38188 20047 38228 20056
rect 37804 19962 37844 20047
rect 37996 19962 38036 20047
rect 38188 19928 38228 19937
rect 38284 19928 38324 20728
rect 38228 19888 38324 19928
rect 38380 20768 38420 20777
rect 38188 19879 38228 19888
rect 38380 19853 38420 20728
rect 38572 20768 38612 21307
rect 38764 20852 38804 21568
rect 39052 21365 39092 21568
rect 39148 21608 39188 21617
rect 39148 21449 39188 21568
rect 39244 21608 39284 21619
rect 39244 21533 39284 21568
rect 39340 21608 39380 21617
rect 39380 21568 39668 21608
rect 39340 21559 39380 21568
rect 39243 21524 39285 21533
rect 39243 21484 39244 21524
rect 39284 21484 39285 21524
rect 39243 21475 39285 21484
rect 39147 21440 39189 21449
rect 39147 21400 39148 21440
rect 39188 21400 39189 21440
rect 39147 21391 39189 21400
rect 39532 21440 39572 21449
rect 39051 21356 39093 21365
rect 39051 21316 39052 21356
rect 39092 21316 39093 21356
rect 39051 21307 39093 21316
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 38764 20812 38996 20852
rect 38572 20719 38612 20728
rect 38764 20684 38804 20693
rect 38668 20644 38764 20684
rect 38476 20600 38516 20609
rect 38668 20600 38708 20644
rect 38764 20635 38804 20644
rect 38516 20560 38708 20600
rect 38476 20551 38516 20560
rect 38956 20516 38996 20812
rect 39148 20768 39188 20777
rect 39532 20768 39572 21400
rect 39188 20728 39572 20768
rect 39148 20719 39188 20728
rect 38860 20476 38996 20516
rect 38572 20096 38612 20105
rect 38860 20096 38900 20476
rect 39628 20189 39668 21568
rect 39916 21449 39956 23668
rect 40011 23120 40053 23129
rect 40011 23080 40012 23120
rect 40052 23080 40053 23120
rect 40011 23071 40053 23080
rect 39915 21440 39957 21449
rect 39915 21400 39916 21440
rect 39956 21400 39957 21440
rect 39915 21391 39957 21400
rect 40012 20768 40052 23071
rect 40108 21533 40148 24331
rect 40396 23717 40436 24340
rect 40492 23792 40532 24751
rect 40684 24641 40724 24726
rect 40588 24632 40628 24641
rect 40588 24464 40628 24592
rect 40683 24632 40725 24641
rect 40683 24592 40684 24632
rect 40724 24592 40725 24632
rect 40683 24583 40725 24592
rect 40780 24464 40820 25096
rect 40876 24809 40916 25096
rect 40875 24800 40917 24809
rect 40875 24760 40876 24800
rect 40916 24760 40917 24800
rect 40875 24751 40917 24760
rect 40876 24632 40916 24641
rect 40876 24473 40916 24592
rect 40971 24632 41013 24641
rect 40971 24592 40972 24632
rect 41012 24592 41013 24632
rect 40971 24583 41013 24592
rect 41068 24632 41108 24643
rect 40972 24498 41012 24583
rect 41068 24557 41108 24592
rect 41067 24548 41109 24557
rect 41067 24508 41068 24548
rect 41108 24508 41109 24548
rect 41067 24499 41109 24508
rect 40588 24424 40820 24464
rect 40875 24464 40917 24473
rect 40875 24424 40876 24464
rect 40916 24424 40917 24464
rect 40875 24415 40917 24424
rect 41164 24305 41204 25852
rect 41356 25472 41396 25481
rect 41260 25432 41356 25472
rect 41163 24296 41205 24305
rect 41163 24256 41164 24296
rect 41204 24256 41205 24296
rect 41163 24247 41205 24256
rect 41164 23969 41204 24247
rect 41163 23960 41205 23969
rect 41163 23920 41164 23960
rect 41204 23920 41205 23960
rect 41163 23911 41205 23920
rect 40780 23836 41108 23876
rect 40492 23743 40532 23752
rect 40684 23792 40724 23801
rect 40780 23792 40820 23836
rect 40724 23752 40820 23792
rect 40684 23743 40724 23752
rect 40395 23708 40437 23717
rect 40395 23668 40396 23708
rect 40436 23668 40437 23708
rect 40395 23659 40437 23668
rect 40588 23708 40628 23717
rect 40588 23624 40628 23668
rect 40875 23708 40917 23717
rect 40875 23668 40876 23708
rect 40916 23668 40917 23708
rect 40875 23659 40917 23668
rect 40588 23584 40820 23624
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 40203 22868 40245 22877
rect 40203 22828 40204 22868
rect 40244 22828 40245 22868
rect 40203 22819 40245 22828
rect 40204 22364 40244 22819
rect 40396 22448 40436 22459
rect 40396 22373 40436 22408
rect 40204 22315 40244 22324
rect 40395 22364 40437 22373
rect 40395 22324 40396 22364
rect 40436 22324 40437 22364
rect 40395 22315 40437 22324
rect 40587 22364 40629 22373
rect 40587 22324 40588 22364
rect 40628 22324 40629 22364
rect 40587 22315 40629 22324
rect 40588 22280 40628 22315
rect 40780 22289 40820 23584
rect 40876 23574 40916 23659
rect 41068 23330 41108 23836
rect 41260 23792 41300 25432
rect 41356 25423 41396 25432
rect 41355 24464 41397 24473
rect 41452 24464 41492 25852
rect 41355 24424 41356 24464
rect 41396 24424 41492 24464
rect 41355 24415 41397 24424
rect 41260 23743 41300 23752
rect 41356 23624 41396 24415
rect 41260 23584 41396 23624
rect 41260 23381 41300 23584
rect 40875 23288 40917 23297
rect 40875 23248 40876 23288
rect 40916 23248 40917 23288
rect 41259 23372 41301 23381
rect 41259 23332 41260 23372
rect 41300 23332 41301 23372
rect 41259 23323 41301 23332
rect 41068 23281 41108 23290
rect 40875 23239 40917 23248
rect 40876 23154 40916 23239
rect 40876 22324 41204 22364
rect 40588 22229 40628 22240
rect 40779 22280 40821 22289
rect 40779 22240 40780 22280
rect 40820 22240 40821 22280
rect 40779 22231 40821 22240
rect 40876 22280 40916 22324
rect 40876 22231 40916 22240
rect 41068 22196 41108 22205
rect 40684 22112 40724 22121
rect 41068 22112 41108 22156
rect 40724 22072 41108 22112
rect 40684 22063 40724 22072
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 41067 21776 41109 21785
rect 41067 21736 41068 21776
rect 41108 21736 41109 21776
rect 41067 21727 41109 21736
rect 41068 21608 41108 21727
rect 41164 21692 41204 22324
rect 41260 21785 41300 23323
rect 41355 23288 41397 23297
rect 41355 23248 41356 23288
rect 41396 23248 41397 23288
rect 41355 23239 41397 23248
rect 41356 23204 41396 23239
rect 41356 23153 41396 23164
rect 41452 23120 41492 23129
rect 41452 23060 41492 23080
rect 41452 23020 41588 23060
rect 41451 22952 41493 22961
rect 41451 22912 41452 22952
rect 41492 22912 41493 22952
rect 41451 22903 41493 22912
rect 41452 22280 41492 22903
rect 41548 22709 41588 23020
rect 41547 22700 41589 22709
rect 41547 22660 41548 22700
rect 41588 22660 41589 22700
rect 41547 22651 41589 22660
rect 41452 22231 41492 22240
rect 41259 21776 41301 21785
rect 41259 21736 41260 21776
rect 41300 21736 41301 21776
rect 41259 21727 41301 21736
rect 41548 21701 41588 22651
rect 41644 22373 41684 26095
rect 42220 25976 42260 26776
rect 42220 25927 42260 25936
rect 41739 25892 41781 25901
rect 41739 25852 41740 25892
rect 41780 25852 41781 25892
rect 41739 25843 41781 25852
rect 41740 23465 41780 25843
rect 42604 25808 42644 30136
rect 42795 30008 42837 30017
rect 42795 29968 42796 30008
rect 42836 29968 42837 30008
rect 42795 29959 42837 29968
rect 42796 27497 42836 29959
rect 42891 29168 42933 29177
rect 42891 29128 42892 29168
rect 42932 29128 42933 29168
rect 42891 29119 42933 29128
rect 42795 27488 42837 27497
rect 42795 27448 42796 27488
rect 42836 27448 42837 27488
rect 42795 27439 42837 27448
rect 42796 26564 42836 27439
rect 42892 26648 42932 29119
rect 43468 28841 43508 30640
rect 43564 29756 43604 29765
rect 43564 29009 43604 29716
rect 43852 29177 43892 31312
rect 43948 31303 43988 31312
rect 43947 31016 43989 31025
rect 43947 30976 43948 31016
rect 43988 30976 43989 31016
rect 43947 30967 43989 30976
rect 43948 30680 43988 30967
rect 44140 30680 44180 30689
rect 43988 30640 44084 30680
rect 43948 30631 43988 30640
rect 43947 30512 43989 30521
rect 43947 30472 43948 30512
rect 43988 30472 43989 30512
rect 43947 30463 43989 30472
rect 43948 30378 43988 30463
rect 44044 30101 44084 30640
rect 44140 30185 44180 30640
rect 44235 30680 44277 30689
rect 44235 30640 44236 30680
rect 44276 30640 44277 30680
rect 44235 30631 44277 30640
rect 44236 30546 44276 30631
rect 44428 30512 44468 30521
rect 44139 30176 44181 30185
rect 44139 30136 44140 30176
rect 44180 30136 44181 30176
rect 44139 30127 44181 30136
rect 44043 30092 44085 30101
rect 44043 30052 44044 30092
rect 44084 30052 44085 30092
rect 44043 30043 44085 30052
rect 43948 29840 43988 29849
rect 44428 29840 44468 30472
rect 44524 30269 44564 32152
rect 45676 32117 45716 32824
rect 45868 32864 45908 33067
rect 45868 32815 45908 32824
rect 45964 32864 46004 32875
rect 45964 32789 46004 32824
rect 45963 32780 46005 32789
rect 45963 32740 45964 32780
rect 46004 32740 46005 32780
rect 45963 32731 46005 32740
rect 45772 32696 45812 32705
rect 45772 32276 45812 32656
rect 45868 32276 45908 32285
rect 45772 32236 45868 32276
rect 45868 32227 45908 32236
rect 46156 32192 46196 33100
rect 46252 32864 46292 32873
rect 46252 32369 46292 32824
rect 46251 32360 46293 32369
rect 46251 32320 46252 32360
rect 46292 32320 46293 32360
rect 46251 32311 46293 32320
rect 46252 32192 46292 32201
rect 46156 32152 46252 32192
rect 46252 32143 46292 32152
rect 45675 32108 45717 32117
rect 45675 32068 45676 32108
rect 45716 32068 45717 32108
rect 45675 32059 45717 32068
rect 45676 31940 45716 31949
rect 45003 31688 45045 31697
rect 45003 31648 45004 31688
rect 45044 31648 45045 31688
rect 45003 31639 45045 31648
rect 45004 30773 45044 31639
rect 45099 30932 45141 30941
rect 45099 30892 45100 30932
rect 45140 30892 45141 30932
rect 45099 30883 45141 30892
rect 45003 30764 45045 30773
rect 45003 30724 45004 30764
rect 45044 30724 45045 30764
rect 45003 30715 45045 30724
rect 44907 30680 44949 30689
rect 44907 30640 44908 30680
rect 44948 30640 44949 30680
rect 44907 30631 44949 30640
rect 45004 30680 45044 30715
rect 44523 30260 44565 30269
rect 44523 30220 44524 30260
rect 44564 30220 44565 30260
rect 44523 30211 44565 30220
rect 44524 29849 44564 30211
rect 44908 30101 44948 30631
rect 45004 30629 45044 30640
rect 45100 30680 45140 30883
rect 45100 30353 45140 30640
rect 45196 30680 45236 30689
rect 45099 30344 45141 30353
rect 45099 30304 45100 30344
rect 45140 30304 45141 30344
rect 45099 30295 45141 30304
rect 44907 30092 44949 30101
rect 44907 30052 44908 30092
rect 44948 30052 44949 30092
rect 44907 30043 44949 30052
rect 43988 29800 44468 29840
rect 44523 29840 44565 29849
rect 44523 29800 44524 29840
rect 44564 29800 44565 29840
rect 43948 29791 43988 29800
rect 44523 29791 44565 29800
rect 44811 29840 44853 29849
rect 44811 29800 44812 29840
rect 44852 29800 44853 29840
rect 44811 29791 44853 29800
rect 44812 29706 44852 29791
rect 43851 29168 43893 29177
rect 43851 29128 43852 29168
rect 43892 29128 43893 29168
rect 43851 29119 43893 29128
rect 45100 29168 45140 29177
rect 45196 29168 45236 30640
rect 45676 30605 45716 31900
rect 46059 31604 46101 31613
rect 46059 31564 46060 31604
rect 46100 31564 46101 31604
rect 46059 31555 46101 31564
rect 46060 30689 46100 31555
rect 46155 31352 46197 31361
rect 46155 31312 46156 31352
rect 46196 31312 46197 31352
rect 46155 31303 46197 31312
rect 45868 30680 45908 30689
rect 45675 30596 45717 30605
rect 45675 30556 45676 30596
rect 45716 30556 45717 30596
rect 45675 30547 45717 30556
rect 45291 30428 45333 30437
rect 45291 30388 45292 30428
rect 45332 30388 45333 30428
rect 45291 30379 45333 30388
rect 45140 29128 45236 29168
rect 45292 29168 45332 30379
rect 45676 29597 45716 30547
rect 45675 29588 45717 29597
rect 45675 29548 45676 29588
rect 45716 29548 45717 29588
rect 45675 29539 45717 29548
rect 45100 29119 45140 29128
rect 45292 29119 45332 29128
rect 45388 29168 45428 29177
rect 43563 29000 43605 29009
rect 43563 28960 43564 29000
rect 43604 28960 43605 29000
rect 43563 28951 43605 28960
rect 44716 29000 44756 29009
rect 43467 28832 43509 28841
rect 43467 28792 43468 28832
rect 43508 28792 43509 28832
rect 43467 28783 43509 28792
rect 44619 28580 44661 28589
rect 44619 28540 44620 28580
rect 44660 28540 44661 28580
rect 44619 28531 44661 28540
rect 44620 28446 44660 28531
rect 43213 28328 43253 28337
rect 43213 27992 43253 28288
rect 43563 28328 43605 28337
rect 44620 28328 44660 28337
rect 43563 28288 43564 28328
rect 43604 28288 43605 28328
rect 43563 28279 43605 28288
rect 44524 28288 44620 28328
rect 43213 27952 43316 27992
rect 43179 27656 43221 27665
rect 43276 27656 43316 27952
rect 43564 27824 43604 28279
rect 44332 28160 44372 28169
rect 44332 27833 44372 28120
rect 43564 27775 43604 27784
rect 44331 27824 44373 27833
rect 44331 27784 44332 27824
rect 44372 27784 44373 27824
rect 44331 27775 44373 27784
rect 43084 27616 43180 27656
rect 43220 27616 43316 27656
rect 42988 26816 43028 26844
rect 43084 26825 43124 27616
rect 43179 27607 43221 27616
rect 43180 27588 43220 27607
rect 44524 27329 44564 28288
rect 44620 28279 44660 28288
rect 44716 28001 44756 28960
rect 45099 29000 45141 29009
rect 45099 28960 45100 29000
rect 45140 28960 45141 29000
rect 45099 28951 45141 28960
rect 45100 28866 45140 28951
rect 45388 28589 45428 29128
rect 45676 29000 45716 29009
rect 45868 29000 45908 30640
rect 46059 30680 46101 30689
rect 46059 30640 46060 30680
rect 46100 30640 46101 30680
rect 46059 30631 46101 30640
rect 46060 30546 46100 30631
rect 45963 30428 46005 30437
rect 45963 30388 45964 30428
rect 46004 30388 46005 30428
rect 45963 30379 46005 30388
rect 45964 30294 46004 30379
rect 46156 30185 46196 31303
rect 46348 30941 46388 33100
rect 46636 33032 46676 33664
rect 46732 33704 46772 33713
rect 46732 33209 46772 33664
rect 46731 33200 46773 33209
rect 46731 33160 46732 33200
rect 46772 33160 46773 33200
rect 46731 33151 46773 33160
rect 46444 32992 46676 33032
rect 46347 30932 46389 30941
rect 46347 30892 46348 30932
rect 46388 30892 46389 30932
rect 46347 30883 46389 30892
rect 46444 30773 46484 32992
rect 46540 32864 46580 32873
rect 46540 32453 46580 32824
rect 46636 32864 46676 32873
rect 46732 32864 46772 33151
rect 46828 33125 46868 34168
rect 46827 33116 46869 33125
rect 46827 33076 46828 33116
rect 46868 33076 46869 33116
rect 46827 33067 46869 33076
rect 46924 33032 46964 33041
rect 46924 32873 46964 32992
rect 46676 32824 46772 32864
rect 46923 32864 46965 32873
rect 46923 32824 46924 32864
rect 46964 32824 46965 32864
rect 46636 32815 46676 32824
rect 46923 32815 46965 32824
rect 47116 32864 47156 32873
rect 46539 32444 46581 32453
rect 46539 32404 46540 32444
rect 46580 32404 46581 32444
rect 46539 32395 46581 32404
rect 46635 32360 46677 32369
rect 46635 32320 46636 32360
rect 46676 32320 46677 32360
rect 47116 32360 47156 32824
rect 47308 32864 47348 32873
rect 47211 32780 47253 32789
rect 47211 32740 47212 32780
rect 47252 32740 47253 32780
rect 47211 32731 47253 32740
rect 47212 32646 47252 32731
rect 47308 32453 47348 32824
rect 47307 32444 47349 32453
rect 47307 32404 47308 32444
rect 47348 32404 47349 32444
rect 47307 32395 47349 32404
rect 47116 32320 47252 32360
rect 46635 32311 46677 32320
rect 46539 32108 46581 32117
rect 46539 32068 46540 32108
rect 46580 32068 46581 32108
rect 46539 32059 46581 32068
rect 46443 30764 46485 30773
rect 46443 30724 46444 30764
rect 46484 30724 46485 30764
rect 46443 30715 46485 30724
rect 46252 30680 46292 30689
rect 46155 30176 46197 30185
rect 46155 30136 46156 30176
rect 46196 30136 46197 30176
rect 46155 30127 46197 30136
rect 45963 30092 46005 30101
rect 45963 30052 45964 30092
rect 46004 30052 46005 30092
rect 45963 30043 46005 30052
rect 45964 29958 46004 30043
rect 46156 29840 46196 30127
rect 46252 30092 46292 30640
rect 46348 30680 46388 30689
rect 46348 30437 46388 30640
rect 46540 30680 46580 32059
rect 46540 30605 46580 30640
rect 46539 30596 46581 30605
rect 46539 30556 46540 30596
rect 46580 30556 46581 30596
rect 46539 30547 46581 30556
rect 46347 30428 46389 30437
rect 46347 30388 46348 30428
rect 46388 30388 46389 30428
rect 46347 30379 46389 30388
rect 46540 30428 46580 30437
rect 46252 30043 46292 30052
rect 45964 29672 46004 29681
rect 45964 29252 46004 29632
rect 46059 29420 46101 29429
rect 46059 29380 46060 29420
rect 46100 29380 46101 29420
rect 46059 29371 46101 29380
rect 45964 29203 46004 29212
rect 46060 29168 46100 29371
rect 46060 29119 46100 29128
rect 45716 28960 45908 29000
rect 45676 28951 45716 28960
rect 45387 28580 45429 28589
rect 45387 28540 45388 28580
rect 45428 28540 45429 28580
rect 45387 28531 45429 28540
rect 46156 28496 46196 29800
rect 46348 29840 46388 29849
rect 46348 29429 46388 29800
rect 46540 29840 46580 30388
rect 46540 29791 46580 29800
rect 46347 29420 46389 29429
rect 46347 29380 46348 29420
rect 46388 29380 46389 29420
rect 46347 29371 46389 29380
rect 46155 28456 46196 28496
rect 46348 29168 46388 29177
rect 46636 29168 46676 32311
rect 47115 32192 47157 32201
rect 47115 32152 47116 32192
rect 47156 32152 47157 32192
rect 47115 32143 47157 32152
rect 47116 32058 47156 32143
rect 47212 31361 47252 32320
rect 47404 32201 47444 34336
rect 48459 34376 48501 34385
rect 48459 34336 48460 34376
rect 48500 34336 48501 34376
rect 48459 34327 48501 34336
rect 49228 34376 49268 34385
rect 48556 34208 48596 34217
rect 48556 33209 48596 34168
rect 49228 34133 49268 34336
rect 49420 34376 49460 34385
rect 49227 34124 49269 34133
rect 49227 34084 49228 34124
rect 49268 34084 49269 34124
rect 49227 34075 49269 34084
rect 48940 33704 48980 33713
rect 48748 33664 48940 33704
rect 48555 33200 48597 33209
rect 48555 33160 48556 33200
rect 48596 33160 48597 33200
rect 48555 33151 48597 33160
rect 47595 33116 47637 33125
rect 47595 33076 47596 33116
rect 47636 33076 47637 33116
rect 47595 33067 47637 33076
rect 47596 32982 47636 33067
rect 48075 33032 48117 33041
rect 48075 32992 48076 33032
rect 48116 32992 48117 33032
rect 48075 32983 48117 32992
rect 48076 32898 48116 32983
rect 47500 32864 47540 32873
rect 47403 32192 47445 32201
rect 47403 32152 47404 32192
rect 47444 32152 47445 32192
rect 47403 32143 47445 32152
rect 47211 31352 47253 31361
rect 47211 31312 47212 31352
rect 47252 31312 47253 31352
rect 47211 31303 47253 31312
rect 47500 30689 47540 32824
rect 47691 32864 47733 32873
rect 47691 32824 47692 32864
rect 47732 32824 47733 32864
rect 47691 32815 47733 32824
rect 48267 32864 48309 32873
rect 48267 32824 48268 32864
rect 48308 32824 48309 32864
rect 48267 32815 48309 32824
rect 47692 32730 47732 32815
rect 48268 32730 48308 32815
rect 48267 32444 48309 32453
rect 48267 32404 48268 32444
rect 48308 32404 48309 32444
rect 48267 32395 48309 32404
rect 48268 32360 48308 32395
rect 48268 32309 48308 32320
rect 48459 32192 48501 32201
rect 48459 32152 48460 32192
rect 48500 32152 48501 32192
rect 48459 32143 48501 32152
rect 48460 32058 48500 32143
rect 48364 31520 48404 31529
rect 48075 31184 48117 31193
rect 48075 31144 48076 31184
rect 48116 31144 48117 31184
rect 48075 31135 48117 31144
rect 48076 30764 48116 31135
rect 48076 30715 48116 30724
rect 47499 30680 47541 30689
rect 47499 30640 47500 30680
rect 47540 30640 47541 30680
rect 48364 30680 48404 31480
rect 48556 31352 48596 33151
rect 48651 33032 48693 33041
rect 48651 32992 48652 33032
rect 48692 32992 48693 33032
rect 48651 32983 48693 32992
rect 48652 32864 48692 32983
rect 48652 32815 48692 32824
rect 48748 32360 48788 33664
rect 48940 33655 48980 33664
rect 49131 33704 49173 33713
rect 49131 33664 49132 33704
rect 49172 33664 49173 33704
rect 49131 33655 49173 33664
rect 49228 33704 49268 33713
rect 49132 33570 49172 33655
rect 48940 33452 48980 33461
rect 48844 33412 48940 33452
rect 48844 32873 48884 33412
rect 48940 33403 48980 33412
rect 49035 33116 49077 33125
rect 49035 33076 49036 33116
rect 49076 33076 49077 33116
rect 49035 33067 49077 33076
rect 48939 33032 48981 33041
rect 48939 32992 48940 33032
rect 48980 32992 48981 33032
rect 48939 32983 48981 32992
rect 48843 32864 48885 32873
rect 48843 32824 48844 32864
rect 48884 32824 48885 32864
rect 48843 32815 48885 32824
rect 48940 32360 48980 32983
rect 48748 32311 48788 32320
rect 48844 32320 48980 32360
rect 48844 32192 48884 32320
rect 49036 32276 49076 33067
rect 48844 32143 48884 32152
rect 48940 32236 49076 32276
rect 48940 32192 48980 32236
rect 48843 31772 48885 31781
rect 48843 31732 48844 31772
rect 48884 31732 48885 31772
rect 48843 31723 48885 31732
rect 48844 31604 48884 31723
rect 48844 31555 48884 31564
rect 48556 31303 48596 31312
rect 48651 31352 48693 31361
rect 48651 31312 48652 31352
rect 48692 31312 48693 31352
rect 48651 31303 48693 31312
rect 48844 31352 48884 31361
rect 48652 31218 48692 31303
rect 48844 31025 48884 31312
rect 48843 31016 48885 31025
rect 48843 30976 48844 31016
rect 48884 30976 48885 31016
rect 48843 30967 48885 30976
rect 48460 30680 48500 30689
rect 48364 30640 48460 30680
rect 47499 30631 47541 30640
rect 48460 30631 48500 30640
rect 47115 30596 47157 30605
rect 47115 30556 47116 30596
rect 47156 30556 47157 30596
rect 47115 30547 47157 30556
rect 47020 30512 47060 30521
rect 46924 30472 47020 30512
rect 46924 29840 46964 30472
rect 47020 30463 47060 30472
rect 46924 29791 46964 29800
rect 46388 29128 46676 29168
rect 45100 28337 45140 28422
rect 45771 28412 45813 28421
rect 45771 28372 45772 28412
rect 45812 28372 45813 28412
rect 45771 28363 45813 28372
rect 44812 28328 44852 28337
rect 44812 28085 44852 28288
rect 44907 28328 44949 28337
rect 44907 28288 44908 28328
rect 44948 28288 44949 28328
rect 44907 28279 44949 28288
rect 45099 28328 45141 28337
rect 45099 28288 45100 28328
rect 45140 28288 45141 28328
rect 45099 28279 45141 28288
rect 45196 28328 45236 28337
rect 44908 28194 44948 28279
rect 45196 28244 45236 28288
rect 45187 28204 45236 28244
rect 45292 28328 45332 28337
rect 45187 28160 45227 28204
rect 45004 28120 45227 28160
rect 44811 28076 44853 28085
rect 44811 28036 44812 28076
rect 44852 28036 44853 28076
rect 44811 28027 44853 28036
rect 44715 27992 44757 28001
rect 44715 27952 44716 27992
rect 44756 27952 44757 27992
rect 44715 27943 44757 27952
rect 44619 27908 44661 27917
rect 44619 27868 44620 27908
rect 44660 27868 44661 27908
rect 44619 27859 44661 27868
rect 44523 27320 44565 27329
rect 44523 27280 44524 27320
rect 44564 27280 44565 27320
rect 44523 27271 44565 27280
rect 44620 27161 44660 27859
rect 44715 27656 44757 27665
rect 44715 27616 44716 27656
rect 44756 27616 44757 27656
rect 44715 27607 44757 27616
rect 44716 27522 44756 27607
rect 45004 27488 45044 28120
rect 45099 27656 45141 27665
rect 45099 27616 45100 27656
rect 45140 27616 45141 27656
rect 45099 27607 45141 27616
rect 44812 27448 45044 27488
rect 44619 27152 44661 27161
rect 44619 27112 44620 27152
rect 44660 27112 44661 27152
rect 44619 27103 44661 27112
rect 43083 26816 43125 26825
rect 43028 26776 43084 26816
rect 43124 26776 43125 26816
rect 42988 26767 43028 26776
rect 43083 26767 43125 26776
rect 43563 26816 43605 26825
rect 43563 26776 43564 26816
rect 43604 26776 43605 26816
rect 43563 26767 43605 26776
rect 42892 26608 43028 26648
rect 42796 26524 42932 26564
rect 42028 25768 42644 25808
rect 41739 23456 41781 23465
rect 41739 23416 41740 23456
rect 41780 23416 41781 23456
rect 41739 23407 41781 23416
rect 41740 23120 41780 23407
rect 41835 23288 41877 23297
rect 41835 23248 41836 23288
rect 41876 23248 41877 23288
rect 41835 23239 41877 23248
rect 41740 23071 41780 23080
rect 41836 22952 41876 23239
rect 42028 23060 42068 25768
rect 42796 25472 42836 25481
rect 42700 25432 42796 25472
rect 42315 24632 42357 24641
rect 42315 24592 42316 24632
rect 42356 24592 42357 24632
rect 42315 24583 42357 24592
rect 42700 24632 42740 25432
rect 42796 25423 42836 25432
rect 42700 24583 42740 24592
rect 42316 24498 42356 24583
rect 42124 23792 42164 23801
rect 42124 23129 42164 23752
rect 42123 23120 42165 23129
rect 42123 23080 42124 23120
rect 42164 23080 42165 23120
rect 42123 23071 42165 23080
rect 41740 22912 41876 22952
rect 41932 23020 42068 23060
rect 41643 22364 41685 22373
rect 41643 22324 41644 22364
rect 41684 22324 41685 22364
rect 41643 22315 41685 22324
rect 41164 21643 41204 21652
rect 41547 21692 41589 21701
rect 41547 21652 41548 21692
rect 41588 21652 41589 21692
rect 41547 21643 41589 21652
rect 40107 21524 40149 21533
rect 40107 21484 40108 21524
rect 40148 21484 40149 21524
rect 40107 21475 40149 21484
rect 40012 20719 40052 20728
rect 40971 20600 41013 20609
rect 40971 20560 40972 20600
rect 41012 20560 41013 20600
rect 40971 20551 41013 20560
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 40972 20189 41012 20551
rect 39627 20180 39669 20189
rect 39627 20140 39628 20180
rect 39668 20140 39669 20180
rect 39627 20131 39669 20140
rect 40971 20180 41013 20189
rect 40971 20140 40972 20180
rect 41012 20140 41013 20180
rect 40971 20131 41013 20140
rect 38612 20056 38900 20096
rect 38572 20047 38612 20056
rect 37611 19844 37653 19853
rect 37611 19804 37612 19844
rect 37652 19804 37653 19844
rect 37611 19795 37653 19804
rect 38379 19844 38421 19853
rect 38379 19804 38380 19844
rect 38420 19804 38421 19844
rect 38379 19795 38421 19804
rect 38667 19844 38709 19853
rect 38667 19804 38668 19844
rect 38708 19804 38709 19844
rect 38667 19795 38709 19804
rect 37612 19710 37652 19795
rect 37515 19508 37557 19517
rect 37515 19468 37516 19508
rect 37556 19468 37557 19508
rect 37515 19459 37557 19468
rect 38284 19424 38324 19433
rect 38324 19384 38612 19424
rect 38284 19375 38324 19384
rect 38187 19256 38229 19265
rect 38187 19216 38188 19256
rect 38228 19216 38229 19256
rect 38187 19207 38229 19216
rect 38380 19256 38420 19265
rect 38188 19122 38228 19207
rect 38380 19013 38420 19216
rect 38572 19256 38612 19384
rect 38572 19207 38612 19216
rect 38668 19256 38708 19795
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 39051 19508 39093 19517
rect 39628 19508 39668 20131
rect 40972 20096 41012 20131
rect 40972 20045 41012 20056
rect 41068 20096 41108 21568
rect 41259 21608 41301 21617
rect 41259 21568 41260 21608
rect 41300 21568 41301 21608
rect 41259 21559 41301 21568
rect 41260 21474 41300 21559
rect 41740 21524 41780 22912
rect 41356 21484 41780 21524
rect 41163 20600 41205 20609
rect 41163 20560 41164 20600
rect 41204 20560 41205 20600
rect 41163 20551 41205 20560
rect 41164 20466 41204 20551
rect 41163 20264 41205 20273
rect 41163 20224 41164 20264
rect 41204 20224 41205 20264
rect 41163 20215 41205 20224
rect 41164 20180 41204 20215
rect 41164 20129 41204 20140
rect 41068 20047 41108 20056
rect 41260 20096 41300 20105
rect 41356 20096 41396 21484
rect 41932 21104 41972 23020
rect 42027 22952 42069 22961
rect 42027 22912 42028 22952
rect 42068 22912 42069 22952
rect 42027 22903 42069 22912
rect 42028 22818 42068 22903
rect 42124 22289 42164 23071
rect 42411 23036 42453 23045
rect 42411 22996 42412 23036
rect 42452 22996 42453 23036
rect 42411 22987 42453 22996
rect 42412 22902 42452 22987
rect 42796 22952 42836 22961
rect 42603 22868 42645 22877
rect 42603 22828 42604 22868
rect 42644 22828 42645 22868
rect 42603 22819 42645 22828
rect 42604 22734 42644 22819
rect 42123 22280 42165 22289
rect 42123 22240 42124 22280
rect 42164 22240 42165 22280
rect 42123 22231 42165 22240
rect 42315 22280 42357 22289
rect 42315 22240 42316 22280
rect 42356 22240 42357 22280
rect 42315 22231 42357 22240
rect 42316 22146 42356 22231
rect 42315 21692 42357 21701
rect 42315 21652 42316 21692
rect 42356 21652 42357 21692
rect 42315 21643 42357 21652
rect 42316 21558 42356 21643
rect 42700 21608 42740 21617
rect 42796 21608 42836 22912
rect 42740 21568 42836 21608
rect 42700 21559 42740 21568
rect 42411 21524 42453 21533
rect 42411 21484 42412 21524
rect 42452 21484 42453 21524
rect 42411 21475 42453 21484
rect 42315 21440 42357 21449
rect 42315 21400 42316 21440
rect 42356 21400 42357 21440
rect 42315 21391 42357 21400
rect 41644 21064 41972 21104
rect 41644 20525 41684 21064
rect 41740 20936 41780 20945
rect 41780 20896 41876 20936
rect 41740 20887 41780 20896
rect 41739 20768 41781 20777
rect 41739 20728 41740 20768
rect 41780 20728 41781 20768
rect 41739 20719 41781 20728
rect 41643 20516 41685 20525
rect 41643 20476 41644 20516
rect 41684 20476 41685 20516
rect 41643 20467 41685 20476
rect 41451 20180 41493 20189
rect 41451 20140 41452 20180
rect 41492 20140 41493 20180
rect 41451 20131 41493 20140
rect 41300 20056 41396 20096
rect 41260 20047 41300 20056
rect 41452 20046 41492 20131
rect 39051 19468 39052 19508
rect 39092 19468 39093 19508
rect 39051 19459 39093 19468
rect 39340 19468 39668 19508
rect 40108 19844 40148 19853
rect 41644 19844 41684 20467
rect 41740 19928 41780 20719
rect 41836 20096 41876 20896
rect 41932 20768 41972 20777
rect 41932 20273 41972 20728
rect 42028 20768 42068 20777
rect 41931 20264 41973 20273
rect 41931 20224 41932 20264
rect 41972 20224 41973 20264
rect 41931 20215 41973 20224
rect 41836 20047 41876 20056
rect 41740 19888 41972 19928
rect 41644 19804 41780 19844
rect 39052 19374 39092 19459
rect 39147 19424 39189 19433
rect 39147 19384 39148 19424
rect 39188 19384 39189 19424
rect 39147 19375 39189 19384
rect 38668 19207 38708 19216
rect 38860 19256 38900 19265
rect 38667 19088 38709 19097
rect 38667 19048 38668 19088
rect 38708 19048 38709 19088
rect 38667 19039 38709 19048
rect 38764 19088 38804 19097
rect 38379 19004 38421 19013
rect 38379 18964 38380 19004
rect 38420 18964 38421 19004
rect 38379 18955 38421 18964
rect 37419 18584 37461 18593
rect 37419 18544 37420 18584
rect 37460 18544 37461 18584
rect 37419 18535 37461 18544
rect 37420 18450 37460 18535
rect 38572 18332 38612 18341
rect 38572 17921 38612 18292
rect 37804 17912 37844 17921
rect 37708 17872 37804 17912
rect 37228 17200 37364 17240
rect 37419 17240 37461 17249
rect 37419 17200 37420 17240
rect 37460 17200 37461 17240
rect 36364 17032 36940 17072
rect 36980 17032 37076 17072
rect 37132 17072 37172 17081
rect 36651 16904 36693 16913
rect 36651 16864 36652 16904
rect 36692 16864 36693 16904
rect 36651 16855 36693 16864
rect 36652 16770 36692 16855
rect 36748 16400 36788 16409
rect 36556 16360 36748 16400
rect 36267 16232 36309 16241
rect 36364 16232 36404 16241
rect 36267 16192 36268 16232
rect 36308 16192 36364 16232
rect 36267 16183 36309 16192
rect 36364 16183 36404 16192
rect 36459 16232 36501 16241
rect 36459 16192 36460 16232
rect 36500 16192 36501 16232
rect 36459 16183 36501 16192
rect 36556 16232 36596 16360
rect 36748 16351 36788 16360
rect 36556 16183 36596 16192
rect 36460 16098 36500 16183
rect 36171 16064 36213 16073
rect 36171 16024 36172 16064
rect 36212 16024 36213 16064
rect 36171 16015 36213 16024
rect 36171 15812 36213 15821
rect 36171 15772 36172 15812
rect 36212 15772 36213 15812
rect 36940 15812 36980 17032
rect 37132 16913 37172 17032
rect 37131 16904 37173 16913
rect 37131 16864 37132 16904
rect 37172 16864 37173 16904
rect 37131 16855 37173 16864
rect 37035 16820 37077 16829
rect 37035 16780 37036 16820
rect 37076 16780 37077 16820
rect 37035 16771 37077 16780
rect 37036 16686 37076 16771
rect 37132 16232 37172 16855
rect 37132 16183 37172 16192
rect 37035 16148 37077 16157
rect 37035 16108 37036 16148
rect 37076 16108 37077 16148
rect 37035 16099 37077 16108
rect 37036 16014 37076 16099
rect 36940 15772 37076 15812
rect 36171 15763 36213 15772
rect 36075 15560 36117 15569
rect 36075 15520 36076 15560
rect 36116 15520 36117 15560
rect 36075 15511 36117 15520
rect 36076 15426 36116 15511
rect 36075 14804 36117 14813
rect 36075 14764 36076 14804
rect 36116 14764 36117 14804
rect 36075 14755 36117 14764
rect 35980 14671 36020 14680
rect 36076 14720 36116 14755
rect 36076 14669 36116 14680
rect 36172 14720 36212 15763
rect 36843 15560 36885 15569
rect 36843 15520 36844 15560
rect 36884 15520 36885 15560
rect 36843 15511 36885 15520
rect 36940 15560 36980 15569
rect 36267 15476 36309 15485
rect 36267 15436 36268 15476
rect 36308 15436 36309 15476
rect 36267 15427 36309 15436
rect 36172 14048 36212 14680
rect 36268 14720 36308 15427
rect 36844 14729 36884 15511
rect 36940 14897 36980 15520
rect 36939 14888 36981 14897
rect 36939 14848 36940 14888
rect 36980 14848 36981 14888
rect 36939 14839 36981 14848
rect 36268 14671 36308 14680
rect 36843 14720 36885 14729
rect 36843 14680 36844 14720
rect 36884 14680 36885 14720
rect 36843 14671 36885 14680
rect 36844 14586 36884 14671
rect 36076 14008 36212 14048
rect 36076 13301 36116 14008
rect 36171 13880 36213 13889
rect 36171 13840 36172 13880
rect 36212 13840 36213 13880
rect 36171 13831 36213 13840
rect 36075 13292 36117 13301
rect 36075 13252 36076 13292
rect 36116 13252 36117 13292
rect 36075 13243 36117 13252
rect 36172 13231 36212 13831
rect 36268 13469 36308 13554
rect 36267 13460 36309 13469
rect 36267 13420 36268 13460
rect 36308 13420 36309 13460
rect 36267 13411 36309 13420
rect 36267 13292 36309 13301
rect 36267 13252 36268 13292
rect 36308 13252 36309 13292
rect 36267 13243 36309 13252
rect 36172 13182 36212 13191
rect 36268 13124 36308 13243
rect 37036 13217 37076 15772
rect 37228 14216 37268 17200
rect 37419 17191 37461 17200
rect 37324 17072 37364 17081
rect 37324 16493 37364 17032
rect 37323 16484 37365 16493
rect 37323 16444 37324 16484
rect 37364 16444 37365 16484
rect 37323 16435 37365 16444
rect 37420 16409 37460 17191
rect 37708 17072 37748 17872
rect 37804 17863 37844 17872
rect 38571 17912 38613 17921
rect 38571 17872 38572 17912
rect 38612 17872 38613 17912
rect 38571 17863 38613 17872
rect 37708 17023 37748 17032
rect 38571 17072 38613 17081
rect 38571 17032 38572 17072
rect 38612 17032 38613 17072
rect 38571 17023 38613 17032
rect 37707 16820 37749 16829
rect 37707 16780 37708 16820
rect 37748 16780 37749 16820
rect 37707 16771 37749 16780
rect 37419 16400 37461 16409
rect 37419 16360 37420 16400
rect 37460 16360 37461 16400
rect 37419 16351 37461 16360
rect 37420 16232 37460 16351
rect 37420 15905 37460 16192
rect 37708 16232 37748 16771
rect 37995 16484 38037 16493
rect 37995 16444 37996 16484
rect 38036 16444 38037 16484
rect 37995 16435 38037 16444
rect 37996 16350 38036 16435
rect 37708 16183 37748 16192
rect 37803 16232 37845 16241
rect 37803 16192 37804 16232
rect 37844 16192 37845 16232
rect 37803 16183 37845 16192
rect 37995 16232 38037 16241
rect 37995 16192 37996 16232
rect 38036 16192 38037 16232
rect 37995 16183 38037 16192
rect 37804 15980 37844 16183
rect 37708 15940 37844 15980
rect 37419 15896 37461 15905
rect 37419 15856 37420 15896
rect 37460 15856 37461 15896
rect 37419 15847 37461 15856
rect 37516 15569 37556 15654
rect 37324 15560 37364 15569
rect 37324 15392 37364 15520
rect 37515 15560 37557 15569
rect 37515 15520 37516 15560
rect 37556 15520 37557 15560
rect 37515 15511 37557 15520
rect 37708 15560 37748 15940
rect 37708 15511 37748 15520
rect 37804 15560 37844 15569
rect 37516 15392 37556 15401
rect 37324 15352 37516 15392
rect 37516 15343 37556 15352
rect 37420 14552 37460 14561
rect 37228 14176 37364 14216
rect 37227 14048 37269 14057
rect 37227 14008 37228 14048
rect 37268 14008 37269 14048
rect 37227 13999 37269 14008
rect 37228 13914 37268 13999
rect 37324 13889 37364 14176
rect 37420 14141 37460 14512
rect 37804 14225 37844 15520
rect 37803 14216 37845 14225
rect 37803 14176 37804 14216
rect 37844 14176 37845 14216
rect 37803 14167 37845 14176
rect 37419 14132 37461 14141
rect 37419 14092 37420 14132
rect 37460 14092 37461 14132
rect 37419 14083 37461 14092
rect 37803 14048 37845 14057
rect 37803 14008 37804 14048
rect 37844 14008 37845 14048
rect 37803 13999 37845 14008
rect 37323 13880 37365 13889
rect 37323 13840 37324 13880
rect 37364 13840 37365 13880
rect 37323 13831 37365 13840
rect 37612 13796 37652 13805
rect 37131 13544 37173 13553
rect 37131 13504 37132 13544
rect 37172 13504 37173 13544
rect 37131 13495 37173 13504
rect 36172 13084 36308 13124
rect 36364 13208 36404 13217
rect 36364 13124 36404 13168
rect 36555 13208 36597 13217
rect 36555 13168 36556 13208
rect 36596 13168 36597 13208
rect 36555 13159 36597 13168
rect 36748 13208 36788 13217
rect 36364 13084 36500 13124
rect 36075 12536 36117 12545
rect 36075 12496 36076 12536
rect 36116 12496 36117 12536
rect 36075 12487 36117 12496
rect 36076 11705 36116 12487
rect 35500 11453 35540 11656
rect 35595 11696 35637 11705
rect 35595 11656 35596 11696
rect 35636 11656 35637 11696
rect 35595 11647 35637 11656
rect 36075 11696 36117 11705
rect 36075 11656 36076 11696
rect 36116 11656 36117 11696
rect 36075 11647 36117 11656
rect 36172 11696 36212 13084
rect 36267 12536 36309 12545
rect 36267 12496 36268 12536
rect 36308 12496 36309 12536
rect 36267 12487 36309 12496
rect 36268 12452 36308 12487
rect 36268 12401 36308 12412
rect 36363 12452 36405 12461
rect 36363 12412 36364 12452
rect 36404 12412 36405 12452
rect 36363 12403 36405 12412
rect 36172 11647 36212 11656
rect 36364 11696 36404 12403
rect 36460 12368 36500 13084
rect 36556 13074 36596 13159
rect 36652 13124 36692 13133
rect 36748 13124 36788 13168
rect 37035 13208 37077 13217
rect 37035 13168 37036 13208
rect 37076 13168 37077 13208
rect 37035 13159 37077 13168
rect 36843 13124 36885 13133
rect 36748 13084 36844 13124
rect 36884 13084 36885 13124
rect 36652 12980 36692 13084
rect 36843 13075 36885 13084
rect 36940 13124 36980 13133
rect 36460 12319 36500 12328
rect 36556 12940 36692 12980
rect 36364 11647 36404 11656
rect 36556 11696 36596 12940
rect 36747 12536 36789 12545
rect 36747 12496 36748 12536
rect 36788 12496 36789 12536
rect 36747 12487 36789 12496
rect 36844 12536 36884 13075
rect 36844 12487 36884 12496
rect 36748 12402 36788 12487
rect 36651 12200 36693 12209
rect 36651 12160 36652 12200
rect 36692 12160 36693 12200
rect 36651 12151 36693 12160
rect 36556 11647 36596 11656
rect 36652 11696 36692 12151
rect 36844 11948 36884 11957
rect 36940 11948 36980 13084
rect 37132 12713 37172 13495
rect 37324 13208 37364 13217
rect 37324 12980 37364 13168
rect 37324 12940 37460 12980
rect 37131 12704 37173 12713
rect 37131 12664 37132 12704
rect 37172 12664 37173 12704
rect 37131 12655 37173 12664
rect 37132 12536 37172 12655
rect 37132 12487 37172 12496
rect 37420 12368 37460 12940
rect 37420 12319 37460 12328
rect 36884 11908 36980 11948
rect 36844 11899 36884 11908
rect 36652 11647 36692 11656
rect 36844 11696 36884 11707
rect 35596 11562 35636 11647
rect 36076 11562 36116 11647
rect 36844 11621 36884 11656
rect 36843 11612 36885 11621
rect 36843 11572 36844 11612
rect 36884 11572 36885 11612
rect 36843 11563 36885 11572
rect 36268 11528 36308 11537
rect 35499 11444 35541 11453
rect 35499 11404 35500 11444
rect 35540 11404 35541 11444
rect 35499 11395 35541 11404
rect 35403 11024 35445 11033
rect 35403 10984 35404 11024
rect 35444 10984 35445 11024
rect 36268 11024 36308 11488
rect 36459 11528 36501 11537
rect 36459 11488 36460 11528
rect 36500 11488 36501 11528
rect 36459 11479 36501 11488
rect 36364 11024 36404 11033
rect 36268 10984 36364 11024
rect 35403 10975 35445 10984
rect 36364 10975 36404 10984
rect 36460 11024 36500 11479
rect 37035 11444 37077 11453
rect 37035 11404 37036 11444
rect 37076 11404 37077 11444
rect 37035 11395 37077 11404
rect 36460 10975 36500 10984
rect 36652 11024 36692 11033
rect 36844 11024 36884 11033
rect 36692 10984 36844 11024
rect 36652 10975 36692 10984
rect 36844 10975 36884 10984
rect 36939 11024 36981 11033
rect 36939 10984 36940 11024
rect 36980 10984 36981 11024
rect 36939 10975 36981 10984
rect 37036 11024 37076 11395
rect 37036 10975 37076 10984
rect 37131 11024 37173 11033
rect 37131 10984 37132 11024
rect 37172 10984 37173 11024
rect 37131 10975 37173 10984
rect 36940 10890 36980 10975
rect 37132 10890 37172 10975
rect 36171 10856 36213 10865
rect 36171 10816 36172 10856
rect 36212 10816 36213 10856
rect 36171 10807 36213 10816
rect 36747 10856 36789 10865
rect 36747 10816 36748 10856
rect 36788 10816 36789 10856
rect 36747 10807 36789 10816
rect 36172 10722 36212 10807
rect 36652 10772 36692 10781
rect 36364 10732 36652 10772
rect 36364 10184 36404 10732
rect 36652 10723 36692 10732
rect 36364 10135 36404 10144
rect 36748 10184 36788 10807
rect 36748 10135 36788 10144
rect 37612 10184 37652 13756
rect 37804 11192 37844 13999
rect 37996 11621 38036 16183
rect 38188 15392 38228 15401
rect 38188 14981 38228 15352
rect 38187 14972 38229 14981
rect 38187 14932 38188 14972
rect 38228 14932 38229 14972
rect 38187 14923 38229 14932
rect 38572 14729 38612 17023
rect 38091 14720 38133 14729
rect 38091 14680 38092 14720
rect 38132 14680 38133 14720
rect 38091 14671 38133 14680
rect 38571 14720 38613 14729
rect 38571 14680 38572 14720
rect 38612 14680 38613 14720
rect 38571 14671 38613 14680
rect 38092 14048 38132 14671
rect 38572 14586 38612 14671
rect 38379 14216 38421 14225
rect 38379 14176 38380 14216
rect 38420 14176 38421 14216
rect 38379 14167 38421 14176
rect 38380 14082 38420 14167
rect 38571 14132 38613 14141
rect 38571 14092 38572 14132
rect 38612 14092 38613 14132
rect 38571 14083 38613 14092
rect 38284 14048 38324 14057
rect 38132 14008 38228 14048
rect 38092 13999 38132 14008
rect 38091 13880 38133 13889
rect 38091 13840 38092 13880
rect 38132 13840 38133 13880
rect 38091 13831 38133 13840
rect 38092 11696 38132 13831
rect 38188 13208 38228 14008
rect 38188 12545 38228 13168
rect 38284 13049 38324 14008
rect 38476 14048 38516 14059
rect 38476 13973 38516 14008
rect 38572 14048 38612 14083
rect 38572 13997 38612 14008
rect 38475 13964 38517 13973
rect 38475 13924 38476 13964
rect 38516 13924 38517 13964
rect 38475 13915 38517 13924
rect 38283 13040 38325 13049
rect 38283 13000 38284 13040
rect 38324 13000 38325 13040
rect 38283 12991 38325 13000
rect 38187 12536 38229 12545
rect 38187 12496 38188 12536
rect 38228 12496 38229 12536
rect 38187 12487 38229 12496
rect 38476 11864 38516 11873
rect 38092 11647 38132 11656
rect 38284 11824 38476 11864
rect 38284 11696 38324 11824
rect 38476 11815 38516 11824
rect 38284 11647 38324 11656
rect 37995 11612 38037 11621
rect 37995 11572 37996 11612
rect 38036 11572 38037 11612
rect 37995 11563 38037 11572
rect 38188 11612 38228 11623
rect 38188 11537 38228 11572
rect 38187 11528 38229 11537
rect 38187 11488 38188 11528
rect 38228 11488 38229 11528
rect 38187 11479 38229 11488
rect 37804 11143 37844 11152
rect 37612 10135 37652 10144
rect 38668 10109 38708 19039
rect 38764 18668 38804 19048
rect 38860 18677 38900 19216
rect 38955 19256 38997 19265
rect 38955 19216 38956 19256
rect 38996 19216 38997 19256
rect 38955 19207 38997 19216
rect 38764 18619 38804 18628
rect 38859 18668 38901 18677
rect 38859 18628 38860 18668
rect 38900 18628 38901 18668
rect 38859 18619 38901 18628
rect 38859 13964 38901 13973
rect 38859 13924 38860 13964
rect 38900 13924 38901 13964
rect 38859 13915 38901 13924
rect 38860 13217 38900 13915
rect 38859 13208 38901 13217
rect 38859 13168 38860 13208
rect 38900 13168 38901 13208
rect 38859 13159 38901 13168
rect 38860 11864 38900 13159
rect 38956 12713 38996 19207
rect 39148 18584 39188 19375
rect 39340 19256 39380 19468
rect 39340 19207 39380 19216
rect 39436 19256 39476 19265
rect 39436 19013 39476 19216
rect 39723 19256 39765 19265
rect 39723 19216 39724 19256
rect 39764 19216 39765 19256
rect 39723 19207 39765 19216
rect 39724 19122 39764 19207
rect 39435 19004 39477 19013
rect 39435 18964 39436 19004
rect 39476 18964 39477 19004
rect 39435 18955 39477 18964
rect 40108 18668 40148 19804
rect 40300 19424 40340 19435
rect 40300 19349 40340 19384
rect 40683 19424 40725 19433
rect 40683 19384 40684 19424
rect 40724 19384 40725 19424
rect 40683 19375 40725 19384
rect 40299 19340 40341 19349
rect 40299 19300 40300 19340
rect 40340 19300 40341 19340
rect 40299 19291 40341 19300
rect 40684 19290 40724 19375
rect 41259 19340 41301 19349
rect 41259 19300 41260 19340
rect 41300 19300 41301 19340
rect 41259 19291 41301 19300
rect 41644 19340 41684 19349
rect 41260 19206 41300 19291
rect 41644 19097 41684 19300
rect 41068 19088 41108 19097
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 40971 18668 41013 18677
rect 40108 18628 40184 18668
rect 39964 18584 40004 18593
rect 39148 18535 39188 18544
rect 39724 18544 39964 18584
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 39724 17081 39764 18544
rect 39964 18535 40004 18544
rect 40144 18416 40184 18628
rect 40971 18628 40972 18668
rect 41012 18628 41013 18668
rect 40971 18619 41013 18628
rect 40012 18376 40184 18416
rect 39819 17744 39861 17753
rect 39819 17704 39820 17744
rect 39860 17704 39861 17744
rect 39819 17695 39861 17704
rect 39820 17610 39860 17695
rect 40012 17165 40052 18376
rect 40203 18248 40245 18257
rect 40203 18208 40204 18248
rect 40244 18208 40245 18248
rect 40203 18199 40245 18208
rect 40204 17744 40244 18199
rect 40204 17695 40244 17704
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 40011 17156 40053 17165
rect 40011 17116 40012 17156
rect 40052 17116 40053 17156
rect 40011 17107 40053 17116
rect 39723 17072 39765 17081
rect 39723 17032 39724 17072
rect 39764 17032 39765 17072
rect 39723 17023 39765 17032
rect 40875 16904 40917 16913
rect 40875 16864 40876 16904
rect 40916 16864 40917 16904
rect 40875 16855 40917 16864
rect 39723 16820 39765 16829
rect 39723 16780 39724 16820
rect 39764 16780 39765 16820
rect 39723 16771 39765 16780
rect 39724 16686 39764 16771
rect 40876 16770 40916 16855
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 39915 16652 39957 16661
rect 39915 16612 39916 16652
rect 39956 16612 39957 16652
rect 39915 16603 39957 16612
rect 39627 16232 39669 16241
rect 39916 16232 39956 16603
rect 39627 16192 39628 16232
rect 39668 16192 39669 16232
rect 39627 16183 39669 16192
rect 39820 16192 39916 16232
rect 39052 15688 39476 15728
rect 39052 15560 39092 15688
rect 39052 15511 39092 15520
rect 39147 15560 39189 15569
rect 39147 15520 39148 15560
rect 39188 15520 39189 15560
rect 39147 15511 39189 15520
rect 39244 15560 39284 15569
rect 39148 15426 39188 15511
rect 39244 15401 39284 15520
rect 39243 15392 39285 15401
rect 39243 15352 39244 15392
rect 39284 15352 39285 15392
rect 39243 15343 39285 15352
rect 39436 15392 39476 15688
rect 39628 15653 39668 16183
rect 39627 15644 39669 15653
rect 39627 15604 39628 15644
rect 39668 15604 39669 15644
rect 39627 15595 39669 15604
rect 39436 15343 39476 15352
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 39435 14972 39477 14981
rect 39435 14932 39436 14972
rect 39476 14932 39477 14972
rect 39435 14923 39477 14932
rect 39436 14720 39476 14923
rect 39436 14671 39476 14680
rect 39628 14645 39668 15595
rect 39724 15560 39764 15569
rect 39627 14636 39669 14645
rect 39627 14596 39628 14636
rect 39668 14596 39669 14636
rect 39627 14587 39669 14596
rect 39724 14468 39764 15520
rect 39820 15560 39860 16192
rect 39916 16183 39956 16192
rect 40107 16232 40149 16241
rect 40107 16192 40108 16232
rect 40148 16192 40149 16232
rect 40107 16183 40149 16192
rect 40684 16232 40724 16241
rect 40724 16192 40916 16232
rect 40684 16183 40724 16192
rect 40012 16148 40052 16157
rect 40012 15989 40052 16108
rect 40108 16098 40148 16183
rect 40300 16148 40340 16157
rect 40204 16108 40300 16148
rect 40011 15980 40053 15989
rect 40011 15940 40012 15980
rect 40052 15940 40053 15980
rect 40011 15931 40053 15940
rect 40011 15812 40053 15821
rect 40011 15772 40012 15812
rect 40052 15772 40053 15812
rect 40011 15763 40053 15772
rect 40012 15560 40052 15763
rect 40204 15728 40244 16108
rect 40300 16099 40340 16108
rect 40779 15980 40821 15989
rect 40779 15940 40780 15980
rect 40820 15940 40821 15980
rect 40779 15931 40821 15940
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 40492 15728 40532 15737
rect 40204 15688 40492 15728
rect 40492 15679 40532 15688
rect 40108 15560 40148 15569
rect 40012 15520 40108 15560
rect 39820 15511 39860 15520
rect 40108 15511 40148 15520
rect 40203 15560 40245 15569
rect 40203 15520 40204 15560
rect 40244 15520 40245 15560
rect 40203 15511 40245 15520
rect 40396 15560 40436 15569
rect 40587 15560 40629 15569
rect 40436 15520 40532 15560
rect 40396 15511 40436 15520
rect 40012 14888 40052 14897
rect 39820 14848 40012 14888
rect 39820 14720 39860 14848
rect 40012 14839 40052 14848
rect 40012 14720 40052 14729
rect 39820 14671 39860 14680
rect 39916 14680 40012 14720
rect 39148 14428 39764 14468
rect 39148 14141 39188 14428
rect 39916 14384 39956 14680
rect 40012 14671 40052 14680
rect 40204 14720 40244 15511
rect 40492 15224 40532 15520
rect 40587 15520 40588 15560
rect 40628 15520 40629 15560
rect 40587 15511 40629 15520
rect 40684 15560 40724 15569
rect 40780 15560 40820 15931
rect 40724 15520 40820 15560
rect 40684 15511 40724 15520
rect 40588 15426 40628 15511
rect 40876 15392 40916 16192
rect 40876 15343 40916 15352
rect 40972 15224 41012 18619
rect 41068 18005 41108 19048
rect 41452 19088 41492 19097
rect 41163 18920 41205 18929
rect 41163 18880 41164 18920
rect 41204 18880 41205 18920
rect 41163 18871 41205 18880
rect 41164 18500 41204 18871
rect 41452 18761 41492 19048
rect 41643 19088 41685 19097
rect 41643 19048 41644 19088
rect 41684 19048 41685 19088
rect 41643 19039 41685 19048
rect 41451 18752 41493 18761
rect 41451 18712 41452 18752
rect 41492 18712 41493 18752
rect 41451 18703 41493 18712
rect 41164 18451 41204 18460
rect 41740 18500 41780 19804
rect 41835 19340 41877 19349
rect 41835 19300 41836 19340
rect 41876 19300 41877 19340
rect 41932 19340 41972 19888
rect 42028 19508 42068 20728
rect 42220 20768 42260 20777
rect 42124 20600 42164 20609
rect 42124 20189 42164 20560
rect 42123 20180 42165 20189
rect 42123 20140 42124 20180
rect 42164 20140 42165 20180
rect 42123 20131 42165 20140
rect 42028 19468 42164 19508
rect 42028 19340 42068 19349
rect 41932 19300 42028 19340
rect 41835 19291 41877 19300
rect 42028 19291 42068 19300
rect 41836 19088 41876 19291
rect 41876 19048 42068 19088
rect 41836 19039 41876 19048
rect 41932 18584 41972 18593
rect 41740 18451 41780 18460
rect 41836 18544 41932 18584
rect 41548 18332 41588 18341
rect 41548 18089 41588 18292
rect 41547 18080 41589 18089
rect 41547 18040 41548 18080
rect 41588 18040 41589 18080
rect 41547 18031 41589 18040
rect 41067 17996 41109 18005
rect 41067 17956 41068 17996
rect 41108 17956 41109 17996
rect 41067 17947 41109 17956
rect 41548 17828 41588 18031
rect 41836 17828 41876 18544
rect 41932 18535 41972 18544
rect 41452 17788 41588 17828
rect 41644 17788 41876 17828
rect 41932 18332 41972 18341
rect 41068 17744 41108 17753
rect 41068 17501 41108 17704
rect 41067 17492 41109 17501
rect 41067 17452 41068 17492
rect 41108 17452 41109 17492
rect 41067 17443 41109 17452
rect 41067 17324 41109 17333
rect 41067 17284 41068 17324
rect 41108 17284 41109 17324
rect 41067 17275 41109 17284
rect 41068 16988 41108 17275
rect 41068 16939 41108 16948
rect 41452 16988 41492 17788
rect 41547 17492 41589 17501
rect 41547 17452 41548 17492
rect 41588 17452 41589 17492
rect 41547 17443 41589 17452
rect 41452 16939 41492 16948
rect 41355 16904 41397 16913
rect 41355 16864 41356 16904
rect 41396 16864 41397 16904
rect 41355 16855 41397 16864
rect 41259 16820 41301 16829
rect 40492 15184 41012 15224
rect 41164 16780 41260 16820
rect 41300 16780 41301 16820
rect 40204 14671 40244 14680
rect 40300 14720 40340 14729
rect 40011 14552 40053 14561
rect 40300 14552 40340 14680
rect 40011 14512 40012 14552
rect 40052 14512 40053 14552
rect 40011 14503 40053 14512
rect 40204 14512 40340 14552
rect 39436 14344 39956 14384
rect 39339 14300 39381 14309
rect 39339 14260 39340 14300
rect 39380 14260 39381 14300
rect 39339 14251 39381 14260
rect 39147 14132 39189 14141
rect 39147 14092 39148 14132
rect 39188 14092 39189 14132
rect 39147 14083 39189 14092
rect 39148 14048 39188 14083
rect 39148 13998 39188 14008
rect 39244 14048 39284 14059
rect 39244 13973 39284 14008
rect 39340 14048 39380 14251
rect 39436 14216 39476 14344
rect 40012 14300 40052 14503
rect 39916 14260 40052 14300
rect 39436 14167 39476 14176
rect 39819 14216 39861 14225
rect 39819 14176 39820 14216
rect 39860 14176 39861 14216
rect 39819 14167 39861 14176
rect 39340 13999 39380 14008
rect 39820 14048 39860 14167
rect 39820 13999 39860 14008
rect 39916 14048 39956 14260
rect 40204 14216 40244 14512
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 41067 14384 41109 14393
rect 41067 14344 41068 14384
rect 41108 14344 41109 14384
rect 41067 14335 41109 14344
rect 40012 14176 40244 14216
rect 40012 14132 40052 14176
rect 40012 14083 40052 14092
rect 39916 13999 39956 14008
rect 40108 14048 40148 14057
rect 39243 13964 39285 13973
rect 39243 13924 39244 13964
rect 39284 13924 39285 13964
rect 39243 13915 39285 13924
rect 40108 13889 40148 14008
rect 40300 14048 40340 14057
rect 40107 13880 40149 13889
rect 40107 13840 40108 13880
rect 40148 13840 40149 13880
rect 40107 13831 40149 13840
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 40300 13469 40340 14008
rect 40684 14048 40724 14057
rect 40299 13460 40341 13469
rect 40299 13420 40300 13460
rect 40340 13420 40341 13460
rect 40299 13411 40341 13420
rect 39532 13376 39572 13385
rect 40684 13376 40724 14008
rect 41068 13973 41108 14335
rect 41164 14309 41204 16780
rect 41259 16771 41301 16780
rect 41260 16686 41300 16771
rect 41260 14720 41300 14729
rect 41163 14300 41205 14309
rect 41163 14260 41164 14300
rect 41204 14260 41205 14300
rect 41163 14251 41205 14260
rect 41260 14225 41300 14680
rect 41356 14720 41396 16855
rect 41548 16232 41588 17443
rect 41644 17240 41684 17788
rect 41932 17753 41972 18292
rect 42028 18173 42068 19048
rect 42124 18845 42164 19468
rect 42220 19256 42260 20728
rect 42220 19207 42260 19216
rect 42316 19256 42356 21391
rect 42412 20777 42452 21475
rect 42892 20852 42932 26524
rect 42988 22877 43028 26608
rect 43564 24632 43604 26767
rect 44139 26648 44181 26657
rect 44139 26608 44140 26648
rect 44180 26608 44372 26648
rect 44139 26599 44181 26608
rect 44140 26514 44180 26599
rect 43852 26144 43892 26153
rect 44236 26144 44276 26153
rect 43852 25649 43892 26104
rect 43948 26104 44236 26144
rect 43851 25640 43893 25649
rect 43851 25600 43852 25640
rect 43892 25600 43893 25640
rect 43851 25591 43893 25600
rect 43852 25472 43892 25481
rect 43948 25472 43988 26104
rect 44236 26095 44276 26104
rect 44043 25640 44085 25649
rect 44043 25600 44044 25640
rect 44084 25600 44085 25640
rect 44043 25591 44085 25600
rect 44044 25556 44084 25591
rect 44332 25565 44372 26608
rect 44812 26060 44852 27448
rect 44907 27320 44949 27329
rect 44907 27280 44908 27320
rect 44948 27280 44949 27320
rect 44907 27271 44949 27280
rect 44908 26069 44948 27271
rect 45100 26144 45140 27607
rect 45100 26095 45140 26104
rect 44716 26020 44852 26060
rect 44907 26060 44949 26069
rect 44907 26020 44908 26060
rect 44948 26020 44949 26060
rect 44044 25505 44084 25516
rect 44331 25556 44373 25565
rect 44331 25516 44332 25556
rect 44372 25516 44373 25556
rect 44331 25507 44373 25516
rect 43892 25432 43988 25472
rect 44235 25472 44277 25481
rect 44235 25432 44236 25472
rect 44276 25432 44277 25472
rect 43852 25423 43892 25432
rect 44235 25423 44277 25432
rect 44044 25304 44084 25313
rect 44236 25304 44276 25423
rect 44332 25313 44372 25398
rect 44619 25388 44661 25397
rect 44619 25348 44620 25388
rect 44660 25348 44661 25388
rect 44619 25339 44661 25348
rect 44084 25264 44180 25304
rect 44044 25255 44084 25264
rect 44140 25136 44180 25264
rect 44236 25255 44276 25264
rect 44331 25304 44373 25313
rect 44331 25264 44332 25304
rect 44372 25264 44373 25304
rect 44331 25255 44373 25264
rect 44620 25304 44660 25339
rect 44524 25136 44564 25145
rect 44140 25096 44524 25136
rect 44524 25087 44564 25096
rect 43564 24583 43604 24592
rect 44427 24632 44469 24641
rect 44620 24632 44660 25264
rect 44427 24592 44428 24632
rect 44468 24592 44469 24632
rect 44427 24583 44469 24592
rect 44524 24592 44660 24632
rect 44716 25304 44756 26020
rect 44907 26011 44949 26020
rect 44811 25892 44853 25901
rect 44811 25852 44812 25892
rect 44852 25852 44853 25892
rect 44811 25843 44853 25852
rect 43275 24548 43317 24557
rect 43275 24508 43276 24548
rect 43316 24508 43317 24548
rect 43275 24499 43317 24508
rect 43276 24044 43316 24499
rect 43755 24464 43797 24473
rect 43755 24424 43756 24464
rect 43796 24424 43797 24464
rect 43755 24415 43797 24424
rect 43276 23995 43316 24004
rect 43276 23624 43316 23635
rect 43276 23549 43316 23584
rect 43275 23540 43317 23549
rect 43275 23500 43276 23540
rect 43316 23500 43317 23540
rect 43275 23491 43317 23500
rect 43756 23297 43796 24415
rect 44235 24380 44277 24389
rect 44235 24340 44236 24380
rect 44276 24340 44277 24380
rect 44235 24331 44277 24340
rect 43851 24296 43893 24305
rect 43851 24256 43852 24296
rect 43892 24256 43893 24296
rect 43851 24247 43893 24256
rect 43755 23288 43797 23297
rect 43755 23248 43756 23288
rect 43796 23248 43797 23288
rect 43755 23239 43797 23248
rect 43852 23060 43892 24247
rect 44043 24212 44085 24221
rect 44043 24172 44044 24212
rect 44084 24172 44085 24212
rect 44043 24163 44085 24172
rect 43947 23792 43989 23801
rect 43947 23752 43948 23792
rect 43988 23752 43989 23792
rect 43947 23743 43989 23752
rect 44044 23792 44084 24163
rect 44139 23960 44181 23969
rect 44139 23920 44140 23960
rect 44180 23920 44181 23960
rect 44139 23911 44181 23920
rect 44044 23743 44084 23752
rect 44140 23792 44180 23911
rect 44140 23743 44180 23752
rect 44236 23792 44276 24331
rect 44331 24212 44373 24221
rect 44331 24172 44332 24212
rect 44372 24172 44373 24212
rect 44331 24163 44373 24172
rect 44236 23743 44276 23752
rect 43948 23658 43988 23743
rect 43852 23020 43988 23060
rect 42987 22868 43029 22877
rect 42987 22828 42988 22868
rect 43028 22828 43029 22868
rect 42987 22819 43029 22828
rect 42988 22373 43028 22819
rect 43179 22784 43221 22793
rect 43084 22744 43180 22784
rect 43220 22744 43221 22784
rect 43084 22457 43124 22744
rect 43179 22735 43221 22744
rect 43180 22716 43220 22735
rect 43467 22700 43509 22709
rect 43467 22660 43468 22700
rect 43508 22660 43509 22700
rect 43467 22651 43509 22660
rect 43468 22541 43508 22651
rect 43467 22532 43509 22541
rect 43467 22492 43468 22532
rect 43508 22492 43509 22532
rect 43467 22483 43509 22492
rect 43083 22448 43125 22457
rect 43083 22408 43084 22448
rect 43124 22408 43125 22448
rect 43083 22399 43125 22408
rect 43468 22398 43508 22483
rect 42987 22364 43029 22373
rect 42987 22324 42988 22364
rect 43028 22324 43029 22364
rect 42987 22315 43029 22324
rect 43563 22280 43605 22289
rect 43563 22240 43564 22280
rect 43604 22240 43605 22280
rect 43563 22231 43605 22240
rect 42987 21860 43029 21869
rect 42987 21820 42988 21860
rect 43028 21820 43029 21860
rect 42987 21811 43029 21820
rect 42892 20803 42932 20812
rect 42411 20768 42453 20777
rect 42411 20728 42412 20768
rect 42452 20728 42453 20768
rect 42411 20719 42453 20728
rect 42316 19207 42356 19216
rect 42412 19256 42452 20719
rect 42700 20096 42740 20105
rect 42700 19265 42740 20056
rect 42891 20012 42933 20021
rect 42891 19972 42892 20012
rect 42932 19972 42933 20012
rect 42891 19963 42933 19972
rect 42412 19207 42452 19216
rect 42507 19256 42549 19265
rect 42507 19216 42508 19256
rect 42548 19216 42549 19256
rect 42507 19207 42549 19216
rect 42699 19256 42741 19265
rect 42892 19256 42932 19963
rect 42699 19216 42700 19256
rect 42740 19216 42741 19256
rect 42699 19207 42741 19216
rect 42796 19216 42892 19256
rect 42508 19088 42548 19207
rect 42508 19048 42740 19088
rect 42123 18836 42165 18845
rect 42123 18796 42124 18836
rect 42164 18796 42165 18836
rect 42123 18787 42165 18796
rect 42603 18668 42645 18677
rect 42603 18628 42604 18668
rect 42644 18628 42645 18668
rect 42603 18619 42645 18628
rect 42124 18584 42164 18593
rect 42027 18164 42069 18173
rect 42027 18124 42028 18164
rect 42068 18124 42069 18164
rect 42027 18115 42069 18124
rect 42027 17996 42069 18005
rect 42027 17956 42028 17996
rect 42068 17956 42069 17996
rect 42027 17947 42069 17956
rect 41931 17744 41973 17753
rect 41931 17704 41932 17744
rect 41972 17704 41973 17744
rect 41931 17695 41973 17704
rect 41644 17191 41684 17200
rect 41740 17072 41780 17081
rect 41740 16829 41780 17032
rect 41836 17072 41876 17081
rect 41836 16913 41876 17032
rect 41932 17072 41972 17083
rect 41932 16997 41972 17032
rect 41931 16988 41973 16997
rect 41931 16948 41932 16988
rect 41972 16948 41973 16988
rect 41931 16939 41973 16948
rect 41835 16904 41877 16913
rect 41835 16864 41836 16904
rect 41876 16864 41877 16904
rect 41835 16855 41877 16864
rect 41739 16820 41781 16829
rect 42028 16820 42068 17947
rect 42124 17753 42164 18544
rect 42220 18584 42260 18593
rect 42412 18584 42452 18593
rect 42220 18425 42260 18544
rect 42316 18544 42412 18584
rect 42219 18416 42261 18425
rect 42219 18376 42220 18416
rect 42260 18376 42261 18416
rect 42219 18367 42261 18376
rect 42316 18005 42356 18544
rect 42412 18535 42452 18544
rect 42604 18584 42644 18619
rect 42604 18533 42644 18544
rect 42700 18584 42740 19048
rect 42796 18761 42836 19216
rect 42892 19207 42932 19216
rect 42891 19088 42933 19097
rect 42891 19048 42892 19088
rect 42932 19048 42933 19088
rect 42891 19039 42933 19048
rect 42795 18752 42837 18761
rect 42795 18712 42796 18752
rect 42836 18712 42837 18752
rect 42795 18703 42837 18712
rect 42892 18752 42932 19039
rect 42892 18703 42932 18712
rect 42700 18535 42740 18544
rect 42411 18416 42453 18425
rect 42411 18376 42412 18416
rect 42452 18376 42453 18416
rect 42411 18367 42453 18376
rect 42412 18282 42452 18367
rect 42796 18332 42836 18703
rect 42508 18292 42836 18332
rect 42892 18332 42932 18341
rect 42315 17996 42357 18005
rect 42315 17956 42316 17996
rect 42356 17956 42357 17996
rect 42315 17947 42357 17956
rect 42123 17744 42165 17753
rect 42123 17704 42124 17744
rect 42164 17704 42165 17744
rect 42123 17695 42165 17704
rect 42220 17576 42260 17585
rect 42124 17536 42220 17576
rect 42124 16997 42164 17536
rect 42220 17527 42260 17536
rect 42508 17408 42548 18292
rect 42892 18257 42932 18292
rect 42891 18248 42933 18257
rect 42891 18208 42892 18248
rect 42932 18208 42933 18248
rect 42988 18248 43028 21811
rect 43564 21608 43604 22231
rect 43564 21559 43604 21568
rect 43468 20852 43508 20861
rect 43084 20600 43124 20609
rect 43084 18509 43124 20560
rect 43276 20600 43316 20609
rect 43468 20600 43508 20812
rect 43659 20852 43701 20861
rect 43659 20812 43660 20852
rect 43700 20812 43701 20852
rect 43659 20803 43701 20812
rect 43660 20718 43700 20803
rect 43948 20684 43988 23020
rect 44139 22952 44181 22961
rect 44139 22912 44140 22952
rect 44180 22912 44181 22952
rect 44139 22903 44181 22912
rect 44140 20852 44180 22903
rect 44332 21449 44372 24163
rect 44428 24044 44468 24583
rect 44524 24221 44564 24592
rect 44716 24548 44756 25264
rect 44812 25304 44852 25843
rect 44812 25255 44852 25264
rect 44620 24508 44756 24548
rect 44908 24632 44948 26011
rect 45292 25397 45332 28288
rect 45388 28328 45428 28337
rect 45580 28328 45620 28337
rect 45428 28288 45580 28328
rect 45388 28279 45428 28288
rect 45580 28279 45620 28288
rect 45772 28328 45812 28363
rect 45868 28337 45908 28422
rect 46155 28412 46195 28456
rect 46252 28412 46292 28421
rect 46155 28372 46196 28412
rect 45772 28277 45812 28288
rect 45867 28328 45909 28337
rect 45867 28288 45868 28328
rect 45908 28288 45909 28328
rect 46156 28328 46196 28372
rect 46252 28328 46292 28372
rect 46156 28288 46292 28328
rect 45867 28279 45909 28288
rect 45676 28160 45716 28169
rect 46060 28160 46100 28171
rect 45716 28120 46004 28160
rect 45676 28111 45716 28120
rect 45483 27992 45525 28001
rect 45483 27952 45484 27992
rect 45524 27952 45525 27992
rect 45483 27943 45525 27952
rect 45675 27992 45717 28001
rect 45675 27952 45676 27992
rect 45716 27952 45717 27992
rect 45675 27943 45717 27952
rect 45484 27656 45524 27943
rect 45580 27656 45620 27665
rect 45484 27616 45580 27656
rect 45580 27607 45620 27616
rect 45388 26816 45428 26825
rect 45388 26153 45428 26776
rect 45387 26144 45429 26153
rect 45387 26104 45388 26144
rect 45428 26104 45429 26144
rect 45387 26095 45429 26104
rect 45291 25388 45333 25397
rect 45291 25348 45292 25388
rect 45332 25348 45333 25388
rect 45291 25339 45333 25348
rect 45003 25304 45045 25313
rect 45003 25264 45004 25304
rect 45044 25264 45045 25304
rect 45003 25255 45045 25264
rect 45004 24800 45044 25255
rect 45291 25220 45333 25229
rect 45291 25180 45292 25220
rect 45332 25180 45333 25220
rect 45291 25171 45333 25180
rect 45004 24751 45044 24760
rect 45100 24632 45140 24641
rect 44523 24212 44565 24221
rect 44523 24172 44524 24212
rect 44564 24172 44565 24212
rect 44523 24163 44565 24172
rect 44428 23995 44468 24004
rect 44620 23969 44660 24508
rect 44908 24473 44948 24592
rect 45004 24592 45100 24632
rect 44907 24464 44949 24473
rect 44907 24424 44908 24464
rect 44948 24424 44949 24464
rect 44907 24415 44949 24424
rect 44715 24380 44757 24389
rect 44715 24340 44716 24380
rect 44756 24340 44757 24380
rect 44715 24331 44757 24340
rect 44716 24246 44756 24331
rect 44619 23960 44661 23969
rect 44524 23920 44620 23960
rect 44660 23920 44661 23960
rect 44427 23792 44469 23801
rect 44427 23752 44428 23792
rect 44468 23752 44469 23792
rect 44427 23743 44469 23752
rect 44428 23658 44468 23743
rect 44524 22952 44564 23920
rect 44619 23911 44661 23920
rect 44619 23792 44661 23801
rect 44619 23752 44620 23792
rect 44660 23752 44661 23792
rect 44619 23743 44661 23752
rect 44716 23792 44756 23801
rect 44620 23658 44660 23743
rect 44619 23288 44661 23297
rect 44619 23248 44620 23288
rect 44660 23248 44661 23288
rect 44619 23239 44661 23248
rect 44716 23288 44756 23752
rect 45004 23381 45044 24592
rect 45100 24583 45140 24592
rect 45196 24632 45236 24641
rect 45099 24464 45141 24473
rect 45099 24424 45100 24464
rect 45140 24424 45141 24464
rect 45099 24415 45141 24424
rect 45100 23792 45140 24415
rect 45196 24389 45236 24592
rect 45195 24380 45237 24389
rect 45195 24340 45196 24380
rect 45236 24340 45237 24380
rect 45195 24331 45237 24340
rect 45100 23465 45140 23752
rect 45099 23456 45141 23465
rect 45099 23416 45100 23456
rect 45140 23416 45141 23456
rect 45099 23407 45141 23416
rect 44811 23372 44853 23381
rect 44811 23332 44812 23372
rect 44852 23332 44853 23372
rect 44811 23323 44853 23332
rect 45003 23372 45045 23381
rect 45003 23332 45004 23372
rect 45044 23332 45045 23372
rect 45003 23323 45045 23332
rect 44716 23239 44756 23248
rect 44620 23120 44660 23239
rect 44620 23071 44660 23080
rect 44812 23120 44852 23323
rect 44812 23071 44852 23080
rect 44908 23120 44948 23129
rect 45100 23120 45140 23407
rect 44524 22912 44660 22952
rect 44331 21440 44373 21449
rect 44331 21400 44332 21440
rect 44372 21400 44373 21440
rect 44331 21391 44373 21400
rect 44140 20803 44180 20812
rect 44620 20777 44660 22912
rect 44908 21860 44948 23080
rect 45012 23080 45140 23120
rect 45012 23060 45052 23080
rect 44716 21820 44948 21860
rect 44716 21776 44756 21820
rect 44716 21727 44756 21736
rect 44619 20768 44661 20777
rect 44619 20728 44620 20768
rect 44660 20728 44661 20768
rect 44619 20719 44661 20728
rect 44812 20768 44852 21820
rect 44908 21617 44948 21820
rect 45004 23020 45052 23060
rect 45292 23045 45332 25171
rect 45483 24380 45525 24389
rect 45483 24340 45484 24380
rect 45524 24340 45525 24380
rect 45483 24331 45525 24340
rect 45387 24044 45429 24053
rect 45387 24004 45388 24044
rect 45428 24004 45429 24044
rect 45387 23995 45429 24004
rect 45388 23792 45428 23995
rect 45388 23120 45428 23752
rect 45484 23792 45524 24331
rect 45484 23743 45524 23752
rect 45580 23129 45620 23214
rect 45484 23120 45524 23129
rect 45388 23080 45484 23120
rect 45484 23071 45524 23080
rect 45579 23120 45621 23129
rect 45579 23080 45580 23120
rect 45620 23080 45621 23120
rect 45579 23071 45621 23080
rect 45676 23120 45716 27943
rect 45964 27740 46004 28120
rect 46060 28085 46100 28120
rect 46059 28076 46101 28085
rect 46059 28036 46060 28076
rect 46100 28036 46101 28076
rect 46059 28027 46101 28036
rect 45964 27691 46004 27700
rect 46252 27656 46292 27665
rect 46348 27656 46388 29128
rect 46636 28337 46676 28422
rect 46443 28328 46485 28337
rect 46443 28288 46444 28328
rect 46484 28288 46485 28328
rect 46443 28279 46485 28288
rect 46635 28328 46677 28337
rect 46635 28288 46636 28328
rect 46676 28288 46677 28328
rect 46635 28279 46677 28288
rect 46828 28328 46868 28337
rect 46292 27616 46388 27656
rect 46252 27607 46292 27616
rect 46059 26396 46101 26405
rect 46059 26356 46060 26396
rect 46100 26356 46101 26396
rect 46059 26347 46101 26356
rect 45963 26144 46005 26153
rect 45963 26104 45964 26144
rect 46004 26104 46005 26144
rect 45963 26095 46005 26104
rect 45964 25304 46004 26095
rect 46060 25817 46100 26347
rect 46348 25985 46388 27616
rect 46444 26312 46484 28279
rect 46731 28244 46773 28253
rect 46731 28204 46732 28244
rect 46772 28204 46773 28244
rect 46731 28195 46773 28204
rect 46635 28160 46677 28169
rect 46635 28120 46636 28160
rect 46676 28120 46677 28160
rect 46635 28111 46677 28120
rect 46636 27740 46676 28111
rect 46732 28110 46772 28195
rect 46731 27992 46773 28001
rect 46731 27952 46732 27992
rect 46772 27952 46773 27992
rect 46731 27943 46773 27952
rect 46636 27691 46676 27700
rect 46540 27656 46580 27667
rect 46540 27581 46580 27616
rect 46539 27572 46581 27581
rect 46539 27532 46540 27572
rect 46580 27532 46581 27572
rect 46539 27523 46581 27532
rect 46732 26984 46772 27943
rect 46828 27488 46868 28288
rect 47116 27656 47156 30547
rect 48844 30521 48884 30967
rect 48843 30512 48885 30521
rect 48843 30472 48844 30512
rect 48884 30472 48885 30512
rect 48843 30463 48885 30472
rect 47787 30176 47829 30185
rect 47787 30136 47788 30176
rect 47828 30136 47829 30176
rect 47787 30127 47829 30136
rect 47788 29849 47828 30127
rect 48940 29933 48980 32152
rect 49036 32147 49076 32156
rect 49036 31865 49076 32107
rect 49131 32108 49173 32117
rect 49131 32068 49132 32108
rect 49172 32068 49173 32108
rect 49131 32059 49173 32068
rect 49035 31856 49077 31865
rect 49035 31816 49036 31856
rect 49076 31816 49077 31856
rect 49035 31807 49077 31816
rect 48939 29924 48981 29933
rect 48939 29884 48940 29924
rect 48980 29884 48981 29924
rect 48939 29875 48981 29884
rect 47787 29840 47829 29849
rect 47787 29800 47788 29840
rect 47828 29800 47829 29840
rect 47787 29791 47829 29800
rect 47788 29706 47828 29791
rect 48940 29672 48980 29681
rect 48940 29429 48980 29632
rect 48939 29420 48981 29429
rect 48939 29380 48940 29420
rect 48980 29380 48981 29420
rect 48939 29371 48981 29380
rect 47596 28496 47636 28505
rect 47500 28456 47596 28496
rect 47307 28244 47349 28253
rect 47307 28204 47308 28244
rect 47348 28204 47349 28244
rect 47307 28195 47349 28204
rect 47020 27616 47116 27656
rect 46924 27488 46964 27497
rect 46828 27448 46924 27488
rect 46924 27439 46964 27448
rect 46636 26944 46772 26984
rect 46540 26312 46580 26321
rect 46444 26272 46540 26312
rect 46540 26263 46580 26272
rect 46444 26144 46484 26155
rect 46444 26069 46484 26104
rect 46636 26144 46676 26944
rect 46827 26816 46869 26825
rect 46827 26776 46828 26816
rect 46868 26776 46869 26816
rect 46827 26767 46869 26776
rect 46828 26682 46868 26767
rect 47020 26237 47060 27616
rect 47116 27607 47156 27616
rect 47308 27656 47348 28195
rect 47403 27740 47445 27749
rect 47403 27700 47404 27740
rect 47444 27700 47445 27740
rect 47403 27691 47445 27700
rect 47308 27607 47348 27616
rect 47404 27656 47444 27691
rect 47404 27605 47444 27616
rect 47116 27404 47156 27413
rect 47116 26816 47156 27364
rect 47116 26767 47156 26776
rect 47307 26816 47349 26825
rect 47307 26776 47308 26816
rect 47348 26776 47349 26816
rect 47307 26767 47349 26776
rect 47500 26816 47540 28456
rect 47596 28447 47636 28456
rect 48843 28160 48885 28169
rect 48843 28120 48844 28160
rect 48884 28120 48885 28160
rect 48843 28111 48885 28120
rect 47595 28076 47637 28085
rect 47595 28036 47596 28076
rect 47636 28036 47637 28076
rect 47595 28027 47637 28036
rect 47596 27656 47636 28027
rect 47691 27740 47733 27749
rect 47691 27700 47692 27740
rect 47732 27700 47733 27740
rect 47691 27691 47733 27700
rect 48844 27740 48884 28111
rect 48844 27691 48884 27700
rect 47596 27607 47636 27616
rect 47692 27606 47732 27691
rect 47788 27656 47828 27667
rect 47788 27581 47828 27616
rect 47979 27656 48021 27665
rect 47979 27616 47980 27656
rect 48020 27616 48021 27656
rect 47979 27607 48021 27616
rect 48651 27656 48693 27665
rect 48651 27616 48652 27656
rect 48692 27616 48693 27656
rect 48651 27607 48693 27616
rect 47787 27572 47829 27581
rect 47787 27532 47788 27572
rect 47828 27532 47829 27572
rect 47787 27523 47829 27532
rect 47980 27522 48020 27607
rect 47500 26767 47540 26776
rect 48364 26816 48404 26825
rect 48652 26816 48692 27607
rect 48404 26776 48692 26816
rect 48364 26767 48404 26776
rect 47019 26228 47061 26237
rect 47019 26188 47020 26228
rect 47060 26188 47061 26228
rect 47019 26179 47061 26188
rect 46443 26060 46485 26069
rect 46443 26020 46444 26060
rect 46484 26020 46485 26060
rect 46443 26011 46485 26020
rect 46347 25976 46389 25985
rect 46347 25936 46348 25976
rect 46388 25936 46389 25976
rect 46347 25927 46389 25936
rect 46251 25892 46293 25901
rect 46251 25852 46252 25892
rect 46292 25852 46293 25892
rect 46251 25843 46293 25852
rect 46539 25892 46581 25901
rect 46539 25852 46540 25892
rect 46580 25852 46581 25892
rect 46539 25843 46581 25852
rect 46059 25808 46101 25817
rect 46059 25768 46060 25808
rect 46100 25768 46101 25808
rect 46059 25759 46101 25768
rect 46252 25758 46292 25843
rect 46347 25472 46389 25481
rect 46347 25432 46348 25472
rect 46388 25432 46389 25472
rect 46347 25423 46389 25432
rect 46252 25305 46292 25313
rect 45964 25255 46004 25264
rect 46156 25304 46292 25305
rect 46156 25265 46252 25304
rect 46156 24464 46196 25265
rect 46251 25264 46252 25265
rect 46252 25255 46292 25264
rect 46348 24557 46388 25423
rect 46444 25313 46484 25398
rect 46443 25304 46485 25313
rect 46443 25264 46444 25304
rect 46484 25264 46485 25304
rect 46443 25255 46485 25264
rect 46540 25136 46580 25843
rect 46636 25724 46676 26104
rect 46732 26144 46772 26153
rect 46732 25901 46772 26104
rect 46731 25892 46773 25901
rect 46731 25852 46732 25892
rect 46772 25852 46773 25892
rect 46731 25843 46773 25852
rect 46636 25684 46964 25724
rect 46732 25304 46772 25313
rect 46732 25145 46772 25264
rect 46924 25304 46964 25684
rect 46924 25255 46964 25264
rect 46828 25220 46868 25229
rect 46731 25136 46773 25145
rect 46444 25096 46580 25136
rect 46636 25096 46732 25136
rect 46772 25096 46773 25136
rect 46444 24716 46484 25096
rect 46444 24667 46484 24676
rect 46540 24632 46580 24641
rect 46636 24632 46676 25096
rect 46731 25087 46773 25096
rect 46828 25061 46868 25180
rect 46827 25052 46869 25061
rect 46827 25012 46828 25052
rect 46868 25012 46869 25052
rect 46827 25003 46869 25012
rect 46580 24592 46676 24632
rect 46827 24632 46869 24641
rect 47020 24632 47060 26179
rect 47308 26144 47348 26767
rect 47212 26104 47348 26144
rect 47787 26144 47829 26153
rect 47787 26104 47788 26144
rect 47828 26104 47829 26144
rect 47212 25388 47252 26104
rect 47787 26095 47829 26104
rect 48652 26144 48692 26776
rect 48843 26228 48885 26237
rect 48843 26188 48844 26228
rect 48884 26188 48885 26228
rect 48843 26179 48885 26188
rect 48652 26095 48692 26104
rect 47788 26010 47828 26095
rect 48844 26094 48884 26179
rect 49132 26153 49172 32059
rect 49228 31781 49268 33664
rect 49420 33140 49460 34336
rect 49515 34376 49557 34385
rect 49515 34336 49516 34376
rect 49556 34336 49557 34376
rect 49515 34327 49557 34336
rect 49516 34242 49556 34327
rect 49324 33100 49460 33140
rect 49227 31772 49269 31781
rect 49227 31732 49228 31772
rect 49268 31732 49269 31772
rect 49227 31723 49269 31732
rect 49324 31361 49364 33100
rect 49516 32864 49556 32873
rect 49612 32864 49652 35176
rect 50476 35216 50516 36007
rect 50955 35972 50997 35981
rect 50955 35932 50956 35972
rect 50996 35932 50997 35972
rect 50955 35923 50997 35932
rect 50956 35838 50996 35923
rect 51244 35888 51284 35897
rect 50764 35720 50804 35729
rect 50476 35167 50516 35176
rect 50668 35680 50764 35720
rect 50475 35048 50517 35057
rect 50475 35008 50476 35048
rect 50516 35008 50517 35048
rect 50475 34999 50517 35008
rect 50379 34712 50421 34721
rect 50379 34672 50380 34712
rect 50420 34672 50421 34712
rect 50379 34663 50421 34672
rect 50091 34124 50133 34133
rect 50091 34084 50092 34124
rect 50132 34084 50133 34124
rect 50091 34075 50133 34084
rect 50092 33140 50132 34075
rect 49556 32824 49652 32864
rect 49516 32815 49556 32824
rect 49420 32192 49460 32203
rect 49612 32201 49652 32824
rect 49804 33100 50132 33140
rect 49420 32117 49460 32152
rect 49611 32192 49653 32201
rect 49611 32152 49612 32192
rect 49652 32152 49653 32192
rect 49611 32143 49653 32152
rect 49419 32108 49461 32117
rect 49419 32068 49420 32108
rect 49460 32068 49461 32108
rect 49419 32059 49461 32068
rect 49612 31940 49652 32143
rect 49515 31520 49557 31529
rect 49515 31480 49516 31520
rect 49556 31480 49557 31520
rect 49515 31471 49557 31480
rect 49228 31352 49268 31361
rect 49228 29849 49268 31312
rect 49323 31352 49365 31361
rect 49323 31312 49324 31352
rect 49364 31312 49365 31352
rect 49323 31303 49365 31312
rect 49420 31352 49460 31361
rect 49323 31184 49365 31193
rect 49323 31144 49324 31184
rect 49364 31144 49365 31184
rect 49323 31135 49365 31144
rect 49324 31050 49364 31135
rect 49420 30857 49460 31312
rect 49516 31352 49556 31471
rect 49516 31303 49556 31312
rect 49419 30848 49461 30857
rect 49419 30808 49420 30848
rect 49460 30808 49461 30848
rect 49419 30799 49461 30808
rect 49324 30680 49364 30689
rect 49612 30680 49652 31900
rect 49708 31529 49748 31614
rect 49707 31520 49749 31529
rect 49707 31480 49708 31520
rect 49748 31480 49749 31520
rect 49707 31471 49749 31480
rect 49708 31352 49748 31361
rect 49804 31352 49844 33100
rect 50091 33032 50133 33041
rect 50091 32992 50092 33032
rect 50132 32992 50133 33032
rect 50091 32983 50133 32992
rect 49995 31772 50037 31781
rect 49995 31732 49996 31772
rect 50036 31732 50037 31772
rect 49995 31723 50037 31732
rect 49748 31312 49844 31352
rect 49708 31303 49748 31312
rect 49364 30640 49652 30680
rect 49324 30269 49364 30640
rect 49419 30512 49461 30521
rect 49419 30472 49420 30512
rect 49460 30472 49461 30512
rect 49419 30463 49461 30472
rect 49323 30260 49365 30269
rect 49323 30220 49324 30260
rect 49364 30220 49365 30260
rect 49323 30211 49365 30220
rect 49324 29924 49364 29933
rect 49227 29840 49269 29849
rect 49227 29800 49228 29840
rect 49268 29800 49269 29840
rect 49227 29791 49269 29800
rect 49324 28664 49364 29884
rect 49420 29084 49460 30463
rect 49804 30008 49844 31312
rect 49900 31352 49940 31361
rect 49900 30773 49940 31312
rect 49996 31352 50036 31723
rect 49996 31303 50036 31312
rect 49899 30764 49941 30773
rect 49899 30724 49900 30764
rect 49940 30724 49941 30764
rect 49899 30715 49941 30724
rect 50092 30008 50132 32983
rect 50284 31352 50324 31361
rect 50380 31352 50420 34663
rect 50476 34385 50516 34999
rect 50475 34376 50517 34385
rect 50475 34336 50476 34376
rect 50516 34336 50517 34376
rect 50475 34327 50517 34336
rect 50572 34376 50612 34385
rect 50476 34242 50516 34327
rect 50572 33125 50612 34336
rect 50668 34376 50708 35680
rect 50764 35671 50804 35680
rect 50860 35216 50900 35225
rect 50860 34628 50900 35176
rect 51052 35048 51092 35057
rect 51244 35048 51284 35848
rect 51435 35888 51477 35897
rect 52396 35888 52436 35897
rect 51435 35848 51436 35888
rect 51476 35848 51477 35888
rect 51435 35839 51477 35848
rect 52204 35848 52396 35888
rect 51340 35804 51380 35813
rect 51340 35384 51380 35764
rect 51436 35754 51476 35839
rect 52012 35804 52052 35813
rect 52052 35764 52148 35804
rect 52012 35755 52052 35764
rect 51340 35344 51572 35384
rect 51340 35216 51380 35225
rect 51340 35057 51380 35176
rect 51435 35216 51477 35225
rect 51435 35176 51436 35216
rect 51476 35176 51477 35216
rect 51435 35167 51477 35176
rect 51436 35082 51476 35167
rect 51532 35141 51572 35344
rect 51627 35300 51669 35309
rect 51627 35260 51628 35300
rect 51668 35260 51669 35300
rect 52108 35300 52148 35764
rect 52204 35384 52244 35848
rect 52396 35839 52436 35848
rect 52779 35888 52821 35897
rect 52779 35848 52780 35888
rect 52820 35848 52821 35888
rect 52779 35839 52821 35848
rect 53260 35877 53300 35886
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 52204 35344 52532 35384
rect 52108 35260 52244 35300
rect 51627 35251 51669 35260
rect 51531 35132 51573 35141
rect 51531 35092 51532 35132
rect 51572 35092 51573 35132
rect 51531 35083 51573 35092
rect 51092 35008 51284 35048
rect 51339 35048 51381 35057
rect 51339 35008 51340 35048
rect 51380 35008 51381 35048
rect 51052 34999 51092 35008
rect 51339 34999 51381 35008
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 51532 34637 51572 35083
rect 50956 34628 50996 34637
rect 50860 34588 50956 34628
rect 50956 34579 50996 34588
rect 51147 34628 51189 34637
rect 51147 34588 51148 34628
rect 51188 34588 51189 34628
rect 51147 34579 51189 34588
rect 51531 34628 51573 34637
rect 51531 34588 51532 34628
rect 51572 34588 51573 34628
rect 51531 34579 51573 34588
rect 50571 33116 50613 33125
rect 50571 33076 50572 33116
rect 50612 33076 50613 33116
rect 50571 33067 50613 33076
rect 50668 33041 50708 34336
rect 50764 34376 50804 34385
rect 50956 34376 50996 34385
rect 50804 34336 50956 34376
rect 50764 34327 50804 34336
rect 50956 34327 50996 34336
rect 51148 34376 51188 34579
rect 51243 34544 51285 34553
rect 51243 34504 51244 34544
rect 51284 34504 51285 34544
rect 51243 34495 51285 34504
rect 51148 34327 51188 34336
rect 51244 34376 51284 34495
rect 51244 34327 51284 34336
rect 51628 34376 51668 35251
rect 51724 35216 51764 35225
rect 52012 35216 52052 35225
rect 51724 34721 51764 35176
rect 51916 35176 52012 35216
rect 51723 34712 51765 34721
rect 51723 34672 51724 34712
rect 51764 34672 51765 34712
rect 51723 34663 51765 34672
rect 51724 34544 51764 34553
rect 51916 34544 51956 35176
rect 52012 35167 52052 35176
rect 52108 35202 52148 35211
rect 52108 35141 52148 35162
rect 52107 35132 52149 35141
rect 52107 35092 52108 35132
rect 52148 35092 52149 35132
rect 52107 35083 52149 35092
rect 52108 35067 52148 35083
rect 52204 34964 52244 35260
rect 52299 35216 52341 35225
rect 52299 35176 52300 35216
rect 52340 35176 52341 35216
rect 52299 35167 52341 35176
rect 52300 35082 52340 35167
rect 52492 35048 52532 35344
rect 52492 34999 52532 35008
rect 52300 34964 52340 34973
rect 52204 34924 52300 34964
rect 52300 34915 52340 34924
rect 52780 34721 52820 35839
rect 53260 35645 53300 35837
rect 54412 35720 54452 35731
rect 54412 35645 54452 35680
rect 53259 35636 53301 35645
rect 53259 35596 53260 35636
rect 53300 35596 53301 35636
rect 53259 35587 53301 35596
rect 54411 35636 54453 35645
rect 54411 35596 54412 35636
rect 54452 35596 54453 35636
rect 54411 35587 54453 35596
rect 54412 35309 54452 35587
rect 55180 35393 55220 35478
rect 55372 35468 55412 37351
rect 55468 36476 55508 37360
rect 55659 37400 55701 37409
rect 55659 37360 55660 37400
rect 55700 37360 55701 37400
rect 55659 37351 55701 37360
rect 55756 37400 55796 37409
rect 55564 37232 55604 37241
rect 55564 36821 55604 37192
rect 55659 37232 55701 37241
rect 55659 37192 55660 37232
rect 55700 37192 55701 37232
rect 55659 37183 55701 37192
rect 55563 36812 55605 36821
rect 55563 36772 55564 36812
rect 55604 36772 55605 36812
rect 55563 36763 55605 36772
rect 55660 36728 55700 37183
rect 55756 36905 55796 37360
rect 55948 37400 55988 37939
rect 55948 37351 55988 37360
rect 56332 37400 56372 37409
rect 56428 37400 56468 38032
rect 57291 38072 57333 38081
rect 57291 38032 57292 38072
rect 57332 38032 57333 38072
rect 57291 38023 57333 38032
rect 57484 37988 57524 37997
rect 56372 37360 56468 37400
rect 57195 37400 57237 37409
rect 57195 37360 57196 37400
rect 57236 37360 57237 37400
rect 56332 37351 56372 37360
rect 57195 37351 57237 37360
rect 57196 37266 57236 37351
rect 57484 37325 57524 37948
rect 57483 37316 57525 37325
rect 57483 37276 57484 37316
rect 57524 37276 57525 37316
rect 57483 37267 57525 37276
rect 56715 37232 56757 37241
rect 56715 37192 56716 37232
rect 56756 37192 56757 37232
rect 56715 37183 56757 37192
rect 55755 36896 55797 36905
rect 55755 36856 55756 36896
rect 55796 36856 55797 36896
rect 55755 36847 55797 36856
rect 55660 36679 55700 36688
rect 56235 36644 56277 36653
rect 56235 36604 56236 36644
rect 56276 36604 56277 36644
rect 56235 36595 56277 36604
rect 55468 36436 55700 36476
rect 55660 36056 55700 36436
rect 55660 36016 55796 36056
rect 55756 35888 55796 36016
rect 55756 35839 55796 35848
rect 55852 35888 55892 35897
rect 55467 35804 55509 35813
rect 55467 35764 55468 35804
rect 55508 35764 55509 35804
rect 55467 35755 55509 35764
rect 55372 35428 55422 35468
rect 55179 35384 55221 35393
rect 55382 35384 55422 35428
rect 55179 35344 55180 35384
rect 55220 35344 55221 35384
rect 55179 35335 55221 35344
rect 55372 35344 55422 35384
rect 54411 35300 54453 35309
rect 54411 35260 54412 35300
rect 54452 35260 54453 35300
rect 54411 35251 54453 35260
rect 54795 35300 54837 35309
rect 54795 35260 54796 35300
rect 54836 35260 54837 35300
rect 54795 35251 54837 35260
rect 55275 35300 55317 35309
rect 55372 35300 55412 35344
rect 55275 35260 55276 35300
rect 55316 35260 55412 35300
rect 55275 35251 55317 35260
rect 54700 35216 54740 35225
rect 52779 34712 52821 34721
rect 52779 34672 52780 34712
rect 52820 34672 52821 34712
rect 52779 34663 52821 34672
rect 52204 34553 52244 34638
rect 51764 34504 51956 34544
rect 52203 34544 52245 34553
rect 52203 34504 52204 34544
rect 52244 34504 52245 34544
rect 51724 34495 51764 34504
rect 52203 34495 52245 34504
rect 52684 34544 52724 34553
rect 52724 34504 52820 34544
rect 52684 34495 52724 34504
rect 51628 34327 51668 34336
rect 51819 34376 51861 34385
rect 51819 34336 51820 34376
rect 51860 34336 51861 34376
rect 51819 34327 51861 34336
rect 52204 34376 52244 34385
rect 50955 33704 50997 33713
rect 50955 33664 50956 33704
rect 50996 33664 50997 33704
rect 50955 33655 50997 33664
rect 50667 33032 50709 33041
rect 50667 32992 50668 33032
rect 50708 32992 50709 33032
rect 50667 32983 50709 32992
rect 50859 32864 50901 32873
rect 50859 32824 50860 32864
rect 50900 32824 50901 32864
rect 50859 32815 50901 32824
rect 50860 32730 50900 32815
rect 50956 32780 50996 33655
rect 51820 33461 51860 34327
rect 52204 34133 52244 34336
rect 52395 34376 52437 34385
rect 52395 34336 52396 34376
rect 52436 34336 52437 34376
rect 52395 34327 52437 34336
rect 52492 34376 52532 34385
rect 52396 34242 52436 34327
rect 52492 34217 52532 34336
rect 52491 34208 52533 34217
rect 52491 34168 52492 34208
rect 52532 34168 52533 34208
rect 52491 34159 52533 34168
rect 52203 34124 52245 34133
rect 52203 34084 52204 34124
rect 52244 34084 52245 34124
rect 52203 34075 52245 34084
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 52203 33788 52245 33797
rect 52203 33748 52204 33788
rect 52244 33748 52245 33788
rect 52203 33739 52245 33748
rect 52204 33654 52244 33739
rect 52588 33704 52628 33713
rect 52780 33704 52820 34504
rect 54124 34385 54164 34470
rect 53932 34376 53972 34385
rect 53643 34208 53685 34217
rect 53643 34168 53644 34208
rect 53684 34168 53685 34208
rect 53643 34159 53685 34168
rect 52628 33664 52820 33704
rect 53452 33704 53492 33713
rect 52588 33655 52628 33664
rect 51531 33452 51573 33461
rect 51531 33412 51532 33452
rect 51572 33412 51573 33452
rect 51531 33403 51573 33412
rect 51819 33452 51861 33461
rect 51819 33412 51820 33452
rect 51860 33412 51861 33452
rect 51819 33403 51861 33412
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 51532 33140 51572 33403
rect 51436 33100 51764 33140
rect 51147 33032 51189 33041
rect 51147 32992 51148 33032
rect 51188 32992 51189 33032
rect 51147 32983 51189 32992
rect 51148 32873 51188 32983
rect 50571 32696 50613 32705
rect 50571 32656 50572 32696
rect 50612 32656 50613 32696
rect 50571 32647 50613 32656
rect 50668 32696 50708 32705
rect 50572 32033 50612 32647
rect 50571 32024 50613 32033
rect 50571 31984 50572 32024
rect 50612 31984 50613 32024
rect 50571 31975 50613 31984
rect 50324 31312 50420 31352
rect 50572 31352 50612 31975
rect 50668 31781 50708 32656
rect 50956 32444 50996 32740
rect 50764 32404 50996 32444
rect 51052 32864 51092 32873
rect 50667 31772 50709 31781
rect 50667 31732 50668 31772
rect 50708 31732 50709 31772
rect 50667 31723 50709 31732
rect 50284 30353 50324 31312
rect 50572 31303 50612 31312
rect 50668 31352 50708 31723
rect 50668 31303 50708 31312
rect 50764 31184 50804 32404
rect 51052 32276 51092 32824
rect 51147 32864 51189 32873
rect 51147 32824 51148 32864
rect 51188 32824 51189 32864
rect 51147 32815 51189 32824
rect 51244 32864 51284 32873
rect 51244 32705 51284 32824
rect 51436 32864 51476 33100
rect 51628 33032 51668 33041
rect 51436 32815 51476 32824
rect 51532 32992 51628 33032
rect 51340 32780 51380 32789
rect 51243 32696 51285 32705
rect 51243 32656 51244 32696
rect 51284 32656 51285 32696
rect 51243 32647 51285 32656
rect 50860 32236 51092 32276
rect 50860 31520 50900 32236
rect 51148 32192 51188 32201
rect 50956 32152 51148 32192
rect 50956 31604 50996 32152
rect 51148 32143 51188 32152
rect 51340 31940 51380 32740
rect 51532 32192 51572 32992
rect 51628 32983 51668 32992
rect 51532 32143 51572 32152
rect 51340 31900 51572 31940
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 51148 31604 51188 31613
rect 50956 31564 51148 31604
rect 51148 31555 51188 31564
rect 50860 31480 50996 31520
rect 50956 31478 50996 31480
rect 50956 31429 50996 31438
rect 51148 31361 51188 31446
rect 51147 31352 51189 31361
rect 51147 31312 51148 31352
rect 51188 31312 51189 31352
rect 51147 31303 51189 31312
rect 51340 31352 51380 31361
rect 51340 31184 51380 31312
rect 51436 31352 51476 31361
rect 51532 31352 51572 31900
rect 51627 31436 51669 31445
rect 51627 31396 51628 31436
rect 51668 31396 51669 31436
rect 51627 31387 51669 31396
rect 51476 31312 51572 31352
rect 51436 31303 51476 31312
rect 51628 31302 51668 31387
rect 50764 31144 51380 31184
rect 50859 30848 50901 30857
rect 50859 30808 50860 30848
rect 50900 30808 50901 30848
rect 50859 30799 50901 30808
rect 50379 30764 50421 30773
rect 50379 30724 50380 30764
rect 50420 30724 50421 30764
rect 50379 30715 50421 30724
rect 50860 30764 50900 30799
rect 51724 30773 51764 33100
rect 51819 32780 51861 32789
rect 51819 32740 51820 32780
rect 51860 32740 51861 32780
rect 51819 32731 51861 32740
rect 51820 31604 51860 32731
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 53452 32201 53492 33664
rect 53644 33629 53684 34159
rect 53643 33620 53685 33629
rect 53643 33580 53644 33620
rect 53684 33580 53685 33620
rect 53643 33571 53685 33580
rect 53644 32864 53684 33571
rect 53739 33116 53781 33125
rect 53739 33076 53740 33116
rect 53780 33076 53781 33116
rect 53739 33067 53781 33076
rect 53644 32815 53684 32824
rect 53740 32864 53780 33067
rect 53740 32815 53780 32824
rect 53835 32864 53877 32873
rect 53835 32824 53836 32864
rect 53876 32824 53877 32864
rect 53835 32815 53877 32824
rect 53932 32864 53972 34336
rect 54123 34376 54165 34385
rect 54123 34336 54124 34376
rect 54164 34336 54165 34376
rect 54123 34327 54165 34336
rect 54220 34376 54260 34385
rect 54028 34208 54068 34217
rect 54028 33797 54068 34168
rect 54123 34124 54165 34133
rect 54123 34084 54124 34124
rect 54164 34084 54165 34124
rect 54123 34075 54165 34084
rect 54027 33788 54069 33797
rect 54027 33748 54028 33788
rect 54068 33748 54069 33788
rect 54027 33739 54069 33748
rect 53932 32815 53972 32824
rect 53836 32730 53876 32815
rect 52395 32192 52437 32201
rect 52395 32152 52396 32192
rect 52436 32152 52437 32192
rect 52395 32143 52437 32152
rect 53451 32192 53493 32201
rect 53451 32152 53452 32192
rect 53492 32152 53493 32192
rect 53451 32143 53493 32152
rect 54124 32192 54164 34075
rect 54220 32360 54260 34336
rect 54603 33956 54645 33965
rect 54603 33916 54604 33956
rect 54644 33916 54645 33956
rect 54603 33907 54645 33916
rect 54604 33629 54644 33907
rect 54603 33620 54645 33629
rect 54603 33580 54604 33620
rect 54644 33580 54645 33620
rect 54603 33571 54645 33580
rect 54604 33486 54644 33571
rect 54315 33284 54357 33293
rect 54315 33244 54316 33284
rect 54356 33244 54357 33284
rect 54315 33235 54357 33244
rect 54220 32311 54260 32320
rect 54124 32143 54164 32152
rect 54316 32192 54356 33235
rect 54603 33116 54645 33125
rect 54603 33076 54604 33116
rect 54644 33076 54645 33116
rect 54603 33067 54645 33076
rect 54604 32360 54644 33067
rect 54700 32537 54740 35176
rect 54796 35166 54836 35251
rect 54892 35216 54932 35225
rect 54892 34880 54932 35176
rect 55083 35216 55125 35225
rect 55276 35216 55316 35251
rect 55468 35216 55508 35755
rect 55852 35729 55892 35848
rect 55948 35888 55988 35897
rect 55851 35720 55893 35729
rect 55851 35680 55852 35720
rect 55892 35680 55893 35720
rect 55851 35671 55893 35680
rect 55852 35468 55892 35671
rect 55660 35428 55892 35468
rect 55563 35300 55605 35309
rect 55563 35260 55564 35300
rect 55604 35260 55605 35300
rect 55563 35251 55605 35260
rect 55083 35176 55084 35216
rect 55124 35176 55220 35216
rect 55083 35167 55125 35176
rect 55084 35082 55124 35167
rect 54892 34840 55124 34880
rect 54987 34712 55029 34721
rect 54987 34672 54988 34712
rect 55028 34672 55029 34712
rect 54987 34663 55029 34672
rect 54988 34376 55028 34663
rect 55084 34628 55124 34840
rect 55180 34805 55220 35176
rect 55276 35166 55316 35176
rect 55390 35205 55508 35216
rect 55430 35176 55508 35205
rect 55564 35166 55604 35251
rect 55390 35156 55430 35165
rect 55179 34796 55221 34805
rect 55179 34756 55180 34796
rect 55220 34756 55221 34796
rect 55179 34747 55221 34756
rect 55564 34628 55604 34637
rect 55084 34588 55564 34628
rect 55564 34579 55604 34588
rect 55084 34385 55124 34416
rect 54988 34327 55028 34336
rect 55083 34376 55125 34385
rect 55083 34336 55084 34376
rect 55124 34336 55125 34376
rect 55083 34327 55125 34336
rect 55180 34376 55220 34385
rect 55220 34336 55412 34376
rect 55180 34327 55220 34336
rect 55084 34292 55124 34327
rect 55084 33881 55124 34252
rect 55275 33956 55317 33965
rect 55275 33916 55276 33956
rect 55316 33916 55317 33956
rect 55275 33907 55317 33916
rect 55083 33872 55125 33881
rect 55083 33832 55084 33872
rect 55124 33832 55125 33872
rect 55083 33823 55125 33832
rect 55276 33788 55316 33907
rect 55276 33739 55316 33748
rect 54892 33704 54932 33713
rect 55180 33704 55220 33713
rect 54795 33452 54837 33461
rect 54795 33412 54796 33452
rect 54836 33412 54837 33452
rect 54795 33403 54837 33412
rect 54796 32864 54836 33403
rect 54892 33377 54932 33664
rect 54988 33664 55180 33704
rect 54891 33368 54933 33377
rect 54891 33328 54892 33368
rect 54932 33328 54933 33368
rect 54891 33319 54933 33328
rect 54699 32528 54741 32537
rect 54699 32488 54700 32528
rect 54740 32488 54741 32528
rect 54699 32479 54741 32488
rect 54796 32360 54836 32824
rect 54891 32864 54933 32873
rect 54891 32824 54892 32864
rect 54932 32824 54933 32864
rect 54891 32815 54933 32824
rect 54988 32864 55028 33664
rect 55180 33655 55220 33664
rect 55275 33536 55317 33545
rect 55275 33496 55276 33536
rect 55316 33496 55317 33536
rect 55372 33536 55412 34336
rect 55564 33536 55604 33545
rect 55372 33496 55564 33536
rect 55275 33487 55317 33496
rect 55564 33487 55604 33496
rect 54892 32730 54932 32815
rect 54988 32621 55028 32824
rect 55179 32864 55221 32873
rect 55179 32824 55180 32864
rect 55220 32824 55221 32864
rect 55179 32815 55221 32824
rect 55276 32864 55316 33487
rect 55371 33368 55413 33377
rect 55371 33328 55372 33368
rect 55412 33328 55413 33368
rect 55371 33319 55413 33328
rect 55276 32815 55316 32824
rect 55180 32730 55220 32815
rect 54987 32612 55029 32621
rect 54987 32572 54988 32612
rect 55028 32572 55029 32612
rect 54987 32563 55029 32572
rect 54604 32320 54740 32360
rect 54796 32320 55028 32360
rect 54316 32143 54356 32152
rect 54412 32192 54452 32203
rect 52396 32058 52436 32143
rect 51820 31555 51860 31564
rect 51915 31436 51957 31445
rect 51915 31396 51916 31436
rect 51956 31396 51957 31436
rect 51915 31387 51957 31396
rect 51820 31184 51860 31193
rect 50283 30344 50325 30353
rect 50283 30304 50284 30344
rect 50324 30304 50325 30344
rect 50283 30295 50325 30304
rect 49612 29968 49844 30008
rect 49900 29968 50132 30008
rect 49515 29924 49557 29933
rect 49515 29884 49516 29924
rect 49556 29884 49557 29924
rect 49515 29875 49557 29884
rect 49516 29672 49556 29875
rect 49516 29623 49556 29632
rect 49612 29336 49652 29968
rect 49900 29924 49940 29968
rect 49804 29884 49940 29924
rect 49707 29840 49749 29849
rect 49707 29800 49708 29840
rect 49748 29800 49749 29840
rect 49707 29791 49749 29800
rect 49804 29840 49844 29884
rect 49995 29840 50037 29849
rect 49804 29791 49844 29800
rect 49900 29819 49940 29828
rect 49708 29706 49748 29791
rect 49995 29800 49996 29840
rect 50036 29800 50037 29840
rect 49995 29791 50037 29800
rect 50284 29840 50324 30295
rect 50284 29791 50324 29800
rect 49900 29765 49940 29779
rect 49899 29756 49941 29765
rect 49899 29716 49900 29756
rect 49940 29716 49941 29756
rect 49899 29707 49941 29716
rect 49900 29684 49940 29707
rect 49996 29706 50036 29791
rect 49652 29296 50228 29336
rect 49612 29287 49652 29296
rect 50188 29168 50228 29296
rect 50188 29119 50228 29128
rect 50380 29168 50420 30715
rect 50763 30680 50805 30689
rect 50763 30640 50764 30680
rect 50804 30640 50805 30680
rect 50763 30631 50805 30640
rect 50764 30546 50804 30631
rect 50476 30428 50516 30437
rect 50763 30428 50805 30437
rect 50516 30388 50708 30428
rect 50476 30379 50516 30388
rect 50668 29849 50708 30388
rect 50763 30388 50764 30428
rect 50804 30388 50805 30428
rect 50763 30379 50805 30388
rect 50475 29840 50517 29849
rect 50475 29800 50476 29840
rect 50516 29800 50517 29840
rect 50475 29791 50517 29800
rect 50572 29840 50612 29849
rect 49996 29084 50036 29093
rect 49460 29044 49652 29084
rect 49420 29035 49460 29044
rect 49324 28624 49460 28664
rect 49324 28496 49364 28505
rect 49228 28456 49324 28496
rect 49228 27656 49268 28456
rect 49324 28447 49364 28456
rect 49228 27607 49268 27616
rect 48939 26144 48981 26153
rect 48939 26104 48940 26144
rect 48980 26104 48981 26144
rect 48939 26095 48981 26104
rect 49131 26144 49173 26153
rect 49131 26104 49132 26144
rect 49172 26104 49173 26144
rect 49131 26095 49173 26104
rect 49228 26144 49268 26153
rect 47403 25976 47445 25985
rect 47403 25936 47404 25976
rect 47444 25936 47445 25976
rect 47403 25927 47445 25936
rect 47404 25842 47444 25927
rect 48364 25892 48404 25901
rect 47212 25348 47348 25388
rect 47116 25220 47156 25229
rect 47116 24893 47156 25180
rect 47115 24884 47157 24893
rect 47115 24844 47116 24884
rect 47156 24844 47157 24884
rect 47115 24835 47157 24844
rect 47308 24809 47348 25348
rect 47500 25304 47540 25313
rect 48364 25304 48404 25852
rect 47540 25264 47636 25304
rect 47500 25255 47540 25264
rect 47499 25052 47541 25061
rect 47499 25012 47500 25052
rect 47540 25012 47541 25052
rect 47499 25003 47541 25012
rect 47307 24800 47349 24809
rect 47307 24760 47308 24800
rect 47348 24760 47349 24800
rect 47307 24751 47349 24760
rect 47116 24632 47156 24641
rect 46827 24592 46828 24632
rect 46868 24592 46869 24632
rect 46540 24583 46580 24592
rect 46827 24583 46869 24592
rect 46924 24592 47116 24632
rect 46347 24548 46389 24557
rect 46347 24508 46348 24548
rect 46388 24508 46389 24548
rect 46347 24499 46389 24508
rect 46828 24498 46868 24583
rect 46156 24415 46196 24424
rect 46924 24221 46964 24592
rect 47116 24583 47156 24592
rect 47211 24632 47253 24641
rect 47211 24592 47212 24632
rect 47252 24592 47253 24632
rect 47211 24583 47253 24592
rect 47308 24632 47348 24643
rect 47116 24464 47156 24473
rect 47212 24464 47252 24583
rect 47308 24557 47348 24592
rect 47404 24632 47444 24641
rect 47500 24632 47540 25003
rect 47444 24592 47540 24632
rect 47404 24583 47444 24592
rect 47307 24548 47349 24557
rect 47307 24508 47308 24548
rect 47348 24508 47349 24548
rect 47307 24499 47349 24508
rect 47156 24424 47252 24464
rect 47596 24464 47636 25264
rect 47116 24415 47156 24424
rect 47596 24415 47636 24424
rect 47115 24296 47157 24305
rect 47115 24256 47116 24296
rect 47156 24256 47157 24296
rect 47115 24247 47157 24256
rect 46251 24212 46293 24221
rect 46251 24172 46252 24212
rect 46292 24172 46293 24212
rect 46251 24163 46293 24172
rect 46923 24212 46965 24221
rect 46923 24172 46924 24212
rect 46964 24172 46965 24212
rect 46923 24163 46965 24172
rect 45772 23960 45812 23969
rect 45772 23792 45812 23920
rect 45964 23792 46004 23801
rect 45772 23752 45964 23792
rect 45964 23743 46004 23752
rect 46059 23792 46101 23801
rect 46059 23752 46060 23792
rect 46100 23752 46101 23792
rect 46059 23743 46101 23752
rect 46156 23792 46196 23801
rect 45868 23129 45908 23214
rect 45676 23060 45716 23080
rect 45867 23120 45909 23129
rect 45867 23080 45868 23120
rect 45908 23080 45909 23120
rect 45867 23071 45909 23080
rect 45964 23120 46004 23129
rect 46060 23120 46100 23743
rect 46156 23633 46196 23752
rect 46155 23624 46197 23633
rect 46155 23584 46156 23624
rect 46196 23584 46197 23624
rect 46155 23575 46197 23584
rect 46156 23129 46196 23214
rect 46004 23080 46100 23120
rect 46155 23120 46197 23129
rect 46252 23120 46292 24163
rect 46924 23960 46964 23969
rect 46828 23920 46924 23960
rect 46539 23372 46581 23381
rect 46539 23332 46540 23372
rect 46580 23332 46581 23372
rect 46539 23323 46581 23332
rect 45964 23071 46004 23080
rect 46155 23071 46156 23120
rect 46196 23080 46292 23120
rect 46444 23120 46484 23129
rect 46196 23071 46197 23080
rect 46156 23060 46196 23069
rect 45291 23036 45333 23045
rect 44907 21608 44949 21617
rect 44907 21568 44908 21608
rect 44948 21568 44949 21608
rect 44907 21559 44949 21568
rect 45004 21608 45044 23020
rect 45291 22996 45292 23036
rect 45332 22996 45333 23036
rect 45676 23020 45812 23060
rect 45291 22987 45333 22996
rect 45004 21559 45044 21568
rect 45100 22280 45140 22289
rect 45003 21440 45045 21449
rect 45003 21400 45004 21440
rect 45044 21400 45045 21440
rect 45003 21391 45045 21400
rect 44812 20719 44852 20728
rect 44907 20768 44949 20777
rect 44907 20728 44908 20768
rect 44948 20728 44949 20768
rect 44907 20719 44949 20728
rect 45004 20768 45044 21391
rect 45004 20719 45044 20728
rect 45100 20768 45140 22240
rect 45292 22280 45332 22289
rect 45196 22112 45236 22121
rect 45196 21701 45236 22072
rect 45292 22037 45332 22240
rect 45387 22280 45429 22289
rect 45387 22240 45388 22280
rect 45428 22240 45429 22280
rect 45387 22231 45429 22240
rect 45580 22280 45620 22289
rect 45388 22146 45428 22231
rect 45291 22028 45333 22037
rect 45291 21988 45292 22028
rect 45332 21988 45333 22028
rect 45291 21979 45333 21988
rect 45580 21953 45620 22240
rect 45772 22280 45812 23020
rect 46156 22868 46196 22877
rect 46444 22868 46484 23080
rect 46196 22828 46484 22868
rect 46156 22819 46196 22828
rect 46155 22700 46197 22709
rect 46155 22660 46156 22700
rect 46196 22660 46197 22700
rect 46155 22651 46197 22660
rect 45772 22231 45812 22240
rect 45676 22196 45716 22205
rect 45579 21944 45621 21953
rect 45579 21904 45580 21944
rect 45620 21904 45621 21944
rect 45579 21895 45621 21904
rect 45195 21692 45237 21701
rect 45195 21652 45196 21692
rect 45236 21652 45237 21692
rect 45195 21643 45237 21652
rect 45292 21608 45332 21619
rect 45292 21533 45332 21568
rect 45387 21608 45429 21617
rect 45387 21568 45388 21608
rect 45428 21568 45429 21608
rect 45387 21559 45429 21568
rect 45291 21524 45333 21533
rect 45291 21484 45292 21524
rect 45332 21484 45333 21524
rect 45291 21475 45333 21484
rect 45388 21474 45428 21559
rect 45676 21524 45716 22156
rect 46059 22028 46101 22037
rect 46059 21988 46060 22028
rect 46100 21988 46101 22028
rect 46059 21979 46101 21988
rect 45964 21608 46004 21617
rect 45868 21568 45964 21608
rect 45676 21484 45812 21524
rect 45675 21356 45717 21365
rect 45675 21316 45676 21356
rect 45716 21316 45717 21356
rect 45675 21307 45717 21316
rect 45676 21222 45716 21307
rect 45483 20852 45525 20861
rect 45483 20812 45484 20852
rect 45524 20812 45525 20852
rect 45483 20803 45525 20812
rect 45100 20719 45140 20728
rect 45484 20768 45524 20803
rect 45676 20777 45716 20862
rect 43948 20644 44276 20684
rect 43852 20600 43892 20609
rect 43468 20560 43852 20600
rect 43276 20021 43316 20560
rect 43275 20012 43317 20021
rect 43275 19972 43276 20012
rect 43316 19972 43317 20012
rect 43275 19963 43317 19972
rect 43275 19844 43317 19853
rect 43275 19804 43276 19844
rect 43316 19804 43317 19844
rect 43275 19795 43317 19804
rect 43276 19349 43316 19795
rect 43564 19424 43604 19433
rect 43275 19340 43317 19349
rect 43275 19300 43276 19340
rect 43316 19300 43317 19340
rect 43275 19291 43317 19300
rect 43276 19256 43316 19291
rect 43180 19229 43220 19238
rect 43276 19206 43316 19216
rect 43180 18929 43220 19189
rect 43179 18920 43221 18929
rect 43179 18880 43180 18920
rect 43220 18880 43221 18920
rect 43179 18871 43221 18880
rect 43467 18752 43509 18761
rect 43467 18712 43468 18752
rect 43508 18712 43509 18752
rect 43467 18703 43509 18712
rect 43083 18500 43125 18509
rect 43083 18460 43084 18500
rect 43124 18460 43125 18500
rect 43083 18451 43125 18460
rect 43084 18366 43124 18451
rect 43275 18416 43317 18425
rect 43275 18376 43276 18416
rect 43316 18376 43317 18416
rect 43275 18367 43317 18376
rect 42988 18208 43124 18248
rect 42891 18199 42933 18208
rect 42892 17996 42932 18199
rect 42220 17368 42548 17408
rect 42604 17956 42932 17996
rect 42220 17072 42260 17368
rect 42604 17324 42644 17956
rect 42700 17837 42740 17868
rect 42699 17828 42741 17837
rect 42699 17788 42700 17828
rect 42740 17788 42741 17828
rect 42699 17779 42741 17788
rect 42220 17023 42260 17032
rect 42412 17284 42644 17324
rect 42700 17744 42740 17779
rect 42123 16988 42165 16997
rect 42123 16948 42124 16988
rect 42164 16948 42165 16988
rect 42123 16939 42165 16948
rect 41739 16780 41740 16820
rect 41780 16780 41781 16820
rect 41739 16771 41781 16780
rect 41932 16780 42068 16820
rect 41588 16192 41684 16232
rect 41548 16183 41588 16192
rect 41644 16073 41684 16192
rect 41643 16064 41685 16073
rect 41643 16024 41644 16064
rect 41684 16024 41685 16064
rect 41643 16015 41685 16024
rect 41452 14729 41492 14814
rect 41356 14477 41396 14680
rect 41451 14720 41493 14729
rect 41451 14680 41452 14720
rect 41492 14680 41493 14720
rect 41451 14671 41493 14680
rect 41548 14552 41588 14561
rect 41452 14512 41548 14552
rect 41355 14468 41397 14477
rect 41355 14428 41356 14468
rect 41396 14428 41397 14468
rect 41355 14419 41397 14428
rect 41355 14300 41397 14309
rect 41355 14260 41356 14300
rect 41396 14260 41397 14300
rect 41355 14251 41397 14260
rect 41259 14216 41301 14225
rect 41259 14176 41260 14216
rect 41300 14176 41301 14216
rect 41259 14167 41301 14176
rect 41067 13964 41109 13973
rect 41067 13924 41068 13964
rect 41108 13924 41109 13964
rect 41067 13915 41109 13924
rect 40780 13376 40820 13385
rect 40684 13336 40780 13376
rect 39339 13124 39381 13133
rect 39339 13084 39340 13124
rect 39380 13084 39381 13124
rect 39339 13075 39381 13084
rect 39340 13040 39380 13075
rect 39340 12989 39380 13000
rect 39532 12980 39572 13336
rect 40780 13327 40820 13336
rect 41068 12980 41108 13915
rect 39436 12940 39572 12980
rect 40780 12940 41108 12980
rect 38955 12704 38997 12713
rect 38955 12664 38956 12704
rect 38996 12664 38997 12704
rect 38955 12655 38997 12664
rect 39052 12536 39092 12545
rect 38956 12496 39052 12536
rect 38956 11948 38996 12496
rect 39052 12487 39092 12496
rect 39436 12536 39476 12940
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 39531 12704 39573 12713
rect 39531 12664 39532 12704
rect 39572 12664 39573 12704
rect 39531 12655 39573 12664
rect 39436 12487 39476 12496
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 39436 11948 39476 11957
rect 38956 11908 39436 11948
rect 39436 11899 39476 11908
rect 38860 11824 38996 11864
rect 38859 11696 38901 11705
rect 38859 11656 38860 11696
rect 38900 11656 38901 11696
rect 38859 11647 38901 11656
rect 38764 11612 38804 11621
rect 38764 11033 38804 11572
rect 38763 11024 38805 11033
rect 38763 10984 38764 11024
rect 38804 10984 38805 11024
rect 38763 10975 38805 10984
rect 38764 10436 38804 10975
rect 38860 10613 38900 11647
rect 38859 10604 38901 10613
rect 38859 10564 38860 10604
rect 38900 10564 38901 10604
rect 38859 10555 38901 10564
rect 38804 10396 38900 10436
rect 38764 10387 38804 10396
rect 38667 10100 38709 10109
rect 38667 10060 38668 10100
rect 38708 10060 38709 10100
rect 38667 10051 38709 10060
rect 29163 9512 29205 9521
rect 29163 9472 29164 9512
rect 29204 9472 29205 9512
rect 38860 9512 38900 10396
rect 38956 10184 38996 11824
rect 39532 11705 39572 12655
rect 40299 12536 40341 12545
rect 40299 12496 40300 12536
rect 40340 12496 40341 12536
rect 40299 12487 40341 12496
rect 40300 12402 40340 12487
rect 39147 11696 39189 11705
rect 39147 11656 39148 11696
rect 39188 11656 39189 11696
rect 39147 11647 39189 11656
rect 39436 11696 39476 11705
rect 39148 11562 39188 11647
rect 39339 11612 39381 11621
rect 39436 11612 39476 11656
rect 39531 11696 39573 11705
rect 39531 11656 39532 11696
rect 39572 11656 39573 11696
rect 39531 11647 39573 11656
rect 39628 11696 39668 11705
rect 39339 11572 39340 11612
rect 39380 11572 39476 11612
rect 39339 11563 39381 11572
rect 39628 11537 39668 11656
rect 39724 11696 39764 11705
rect 39627 11528 39669 11537
rect 39627 11488 39628 11528
rect 39668 11488 39669 11528
rect 39627 11479 39669 11488
rect 39435 11024 39477 11033
rect 39435 10984 39436 11024
rect 39476 10984 39477 11024
rect 39435 10975 39477 10984
rect 39436 10890 39476 10975
rect 39724 10688 39764 11656
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 39628 10648 39764 10688
rect 39820 10856 39860 10865
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 39628 10436 39668 10648
rect 38956 10135 38996 10144
rect 39052 10396 39668 10436
rect 39052 10100 39092 10396
rect 39147 10268 39189 10277
rect 39147 10228 39148 10268
rect 39188 10228 39189 10268
rect 39147 10219 39189 10228
rect 39148 10184 39188 10219
rect 39148 10133 39188 10144
rect 39724 10184 39764 10193
rect 39820 10184 39860 10816
rect 40011 10772 40053 10781
rect 40011 10732 40012 10772
rect 40052 10732 40053 10772
rect 40011 10723 40053 10732
rect 39764 10144 39860 10184
rect 39724 10135 39764 10144
rect 39052 10051 39092 10060
rect 39243 10100 39285 10109
rect 39243 10060 39244 10100
rect 39284 10060 39285 10100
rect 39243 10051 39285 10060
rect 39340 10100 39380 10109
rect 39148 9512 39188 9521
rect 38860 9472 39148 9512
rect 29163 9463 29205 9472
rect 39148 9463 39188 9472
rect 39244 9512 39284 10051
rect 39340 9689 39380 10060
rect 39339 9680 39381 9689
rect 39339 9640 39340 9680
rect 39380 9640 39381 9680
rect 39339 9631 39381 9640
rect 39436 9521 39476 9606
rect 39244 9463 39284 9472
rect 39435 9512 39477 9521
rect 39435 9472 39436 9512
rect 39476 9472 39477 9512
rect 39435 9463 39477 9472
rect 39916 9512 39956 9521
rect 39436 9344 39476 9353
rect 39916 9344 39956 9472
rect 40012 9512 40052 10723
rect 40588 10184 40628 10193
rect 40588 10025 40628 10144
rect 40587 10016 40629 10025
rect 40587 9976 40588 10016
rect 40628 9976 40629 10016
rect 40587 9967 40629 9976
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 40780 9689 40820 12940
rect 40875 10100 40917 10109
rect 40875 10060 40876 10100
rect 40916 10060 40917 10100
rect 40875 10051 40917 10060
rect 40107 9680 40149 9689
rect 40107 9640 40108 9680
rect 40148 9640 40149 9680
rect 40107 9631 40149 9640
rect 40779 9680 40821 9689
rect 40779 9640 40780 9680
rect 40820 9640 40821 9680
rect 40779 9631 40821 9640
rect 40108 9546 40148 9631
rect 40683 9596 40725 9605
rect 40683 9556 40684 9596
rect 40724 9556 40725 9596
rect 40683 9547 40725 9556
rect 40012 9463 40052 9472
rect 40203 9512 40245 9521
rect 40203 9472 40204 9512
rect 40244 9472 40245 9512
rect 40203 9463 40245 9472
rect 40587 9512 40629 9521
rect 40587 9472 40588 9512
rect 40628 9472 40629 9512
rect 40587 9463 40629 9472
rect 40684 9512 40724 9547
rect 40204 9378 40244 9463
rect 40588 9378 40628 9463
rect 40684 9461 40724 9472
rect 40780 9512 40820 9631
rect 40780 9463 40820 9472
rect 40876 9512 40916 10051
rect 41356 9605 41396 14251
rect 41452 13208 41492 14512
rect 41548 14503 41588 14512
rect 41548 14048 41588 14057
rect 41644 14048 41684 16015
rect 41836 15560 41876 15569
rect 41932 15560 41972 16780
rect 42027 15644 42069 15653
rect 42027 15604 42028 15644
rect 42068 15604 42069 15644
rect 42027 15595 42069 15604
rect 41876 15520 41972 15560
rect 41836 15511 41876 15520
rect 41588 14008 41684 14048
rect 41836 15308 41876 15317
rect 41548 13999 41588 14008
rect 41547 13460 41589 13469
rect 41547 13420 41548 13460
rect 41588 13420 41589 13460
rect 41547 13411 41589 13420
rect 41548 13326 41588 13411
rect 41548 13208 41588 13217
rect 41452 13168 41548 13208
rect 41548 13159 41588 13168
rect 41739 13208 41781 13217
rect 41739 13168 41740 13208
rect 41780 13168 41781 13208
rect 41739 13159 41781 13168
rect 41836 13208 41876 15268
rect 41932 13889 41972 15520
rect 42028 15560 42068 15595
rect 42028 15509 42068 15520
rect 42124 15560 42164 16939
rect 42219 15644 42261 15653
rect 42219 15604 42220 15644
rect 42260 15604 42261 15644
rect 42219 15595 42261 15604
rect 42124 15511 42164 15520
rect 42027 14720 42069 14729
rect 42027 14680 42028 14720
rect 42068 14680 42069 14720
rect 42027 14671 42069 14680
rect 41931 13880 41973 13889
rect 41931 13840 41932 13880
rect 41972 13840 41973 13880
rect 41931 13831 41973 13840
rect 41836 13159 41876 13168
rect 41740 13074 41780 13159
rect 41452 12704 41492 12715
rect 41452 12629 41492 12664
rect 41451 12620 41493 12629
rect 41451 12580 41452 12620
rect 41492 12580 41493 12620
rect 41451 12571 41493 12580
rect 41452 11789 41492 12571
rect 41739 12536 41781 12545
rect 41739 12496 41740 12536
rect 41780 12496 41781 12536
rect 41739 12487 41781 12496
rect 41451 11780 41493 11789
rect 41451 11740 41452 11780
rect 41492 11740 41493 11780
rect 41451 11731 41493 11740
rect 41548 11024 41588 11033
rect 41740 11024 41780 12487
rect 41835 12284 41877 12293
rect 41835 12244 41836 12284
rect 41876 12244 41877 12284
rect 41835 12235 41877 12244
rect 41836 11696 41876 12235
rect 41836 11647 41876 11656
rect 41932 11696 41972 11705
rect 42028 11696 42068 14671
rect 42220 12536 42260 15595
rect 42315 13880 42357 13889
rect 42315 13840 42316 13880
rect 42356 13840 42357 13880
rect 42315 13831 42357 13840
rect 42316 12881 42356 13831
rect 42412 12980 42452 17284
rect 42508 17072 42548 17081
rect 42508 16241 42548 17032
rect 42604 17072 42644 17083
rect 42604 16997 42644 17032
rect 42603 16988 42645 16997
rect 42603 16948 42604 16988
rect 42644 16948 42645 16988
rect 42603 16939 42645 16948
rect 42700 16820 42740 17704
rect 42891 17744 42933 17753
rect 42891 17704 42892 17744
rect 42932 17704 42933 17744
rect 42891 17695 42933 17704
rect 42988 17744 43028 17753
rect 42795 17660 42837 17669
rect 42795 17620 42796 17660
rect 42836 17620 42837 17660
rect 42795 17611 42837 17620
rect 42796 17526 42836 17611
rect 42892 17610 42932 17695
rect 42891 16904 42933 16913
rect 42891 16864 42892 16904
rect 42932 16864 42933 16904
rect 42891 16855 42933 16864
rect 42604 16780 42740 16820
rect 42507 16232 42549 16241
rect 42507 16192 42508 16232
rect 42548 16192 42549 16232
rect 42507 16183 42549 16192
rect 42604 14729 42644 16780
rect 42892 16770 42932 16855
rect 42699 16652 42741 16661
rect 42699 16612 42700 16652
rect 42740 16612 42741 16652
rect 42699 16603 42741 16612
rect 42700 16484 42740 16603
rect 42700 16435 42740 16444
rect 42988 16484 43028 17704
rect 43084 16988 43124 18208
rect 43179 17660 43221 17669
rect 43179 17620 43180 17660
rect 43220 17620 43221 17660
rect 43179 17611 43221 17620
rect 43180 17526 43220 17611
rect 43276 16988 43316 18367
rect 43371 17324 43413 17333
rect 43371 17284 43372 17324
rect 43412 17284 43413 17324
rect 43371 17275 43413 17284
rect 43084 16939 43124 16948
rect 43180 16948 43316 16988
rect 43180 16820 43220 16948
rect 42988 16435 43028 16444
rect 43084 16780 43220 16820
rect 43276 16820 43316 16829
rect 43372 16820 43412 17275
rect 43316 16780 43412 16820
rect 42891 16232 42933 16241
rect 42891 16192 42892 16232
rect 42932 16192 42933 16232
rect 42891 16183 42933 16192
rect 43084 16232 43124 16780
rect 43276 16771 43316 16780
rect 42892 16098 42932 16183
rect 43084 15653 43124 16192
rect 43276 16148 43316 16157
rect 43276 15905 43316 16108
rect 43275 15896 43317 15905
rect 43275 15856 43276 15896
rect 43316 15856 43317 15896
rect 43275 15847 43317 15856
rect 43083 15644 43125 15653
rect 43083 15604 43084 15644
rect 43124 15604 43125 15644
rect 43083 15595 43125 15604
rect 43084 14888 43124 15595
rect 43468 15224 43508 18703
rect 43564 18584 43604 19384
rect 43660 19004 43700 20560
rect 43852 20551 43892 20560
rect 44236 20012 44276 20644
rect 44908 20634 44948 20719
rect 45484 20717 45524 20728
rect 45675 20768 45717 20777
rect 45675 20728 45676 20768
rect 45716 20728 45717 20768
rect 45675 20719 45717 20728
rect 45772 20768 45812 21484
rect 45772 20719 45812 20728
rect 44332 20600 44372 20609
rect 45580 20600 45620 20609
rect 45868 20600 45908 21568
rect 45964 21559 46004 21568
rect 45963 21356 46005 21365
rect 45963 21316 45964 21356
rect 46004 21316 46005 21356
rect 45963 21307 46005 21316
rect 45964 20768 46004 21307
rect 46060 21020 46100 21979
rect 46060 20777 46100 20980
rect 45964 20719 46004 20728
rect 46059 20768 46101 20777
rect 46059 20728 46060 20768
rect 46100 20728 46101 20768
rect 46059 20719 46101 20728
rect 46156 20768 46196 22651
rect 46444 22448 46484 22457
rect 46251 22280 46293 22289
rect 46251 22240 46252 22280
rect 46292 22240 46293 22280
rect 46251 22231 46293 22240
rect 46252 21020 46292 22231
rect 46348 21608 46388 21617
rect 46444 21608 46484 22408
rect 46388 21568 46484 21608
rect 46348 21559 46388 21568
rect 46348 21020 46388 21029
rect 46252 20980 46348 21020
rect 46348 20971 46388 20980
rect 46156 20719 46196 20728
rect 46347 20768 46389 20777
rect 46347 20728 46348 20768
rect 46388 20728 46389 20768
rect 46347 20719 46389 20728
rect 46540 20768 46580 23323
rect 46731 23204 46773 23213
rect 46731 23164 46732 23204
rect 46772 23164 46773 23204
rect 46731 23155 46773 23164
rect 46635 22280 46677 22289
rect 46635 22240 46636 22280
rect 46676 22240 46677 22280
rect 46635 22231 46677 22240
rect 46540 20719 46580 20728
rect 46636 20768 46676 22231
rect 46732 20777 46772 23155
rect 46828 23120 46868 23920
rect 46924 23911 46964 23920
rect 46828 23071 46868 23080
rect 47116 23060 47156 24247
rect 48364 23969 48404 25264
rect 48460 24464 48500 24473
rect 47691 23960 47733 23969
rect 47691 23920 47692 23960
rect 47732 23920 47733 23960
rect 47691 23911 47733 23920
rect 48363 23960 48405 23969
rect 48363 23920 48364 23960
rect 48404 23920 48405 23960
rect 48363 23911 48405 23920
rect 47692 23120 47732 23911
rect 48364 23792 48404 23801
rect 48460 23792 48500 24424
rect 48555 24296 48597 24305
rect 48555 24256 48556 24296
rect 48596 24256 48597 24296
rect 48555 24247 48597 24256
rect 48404 23752 48500 23792
rect 48364 23743 48404 23752
rect 47980 23708 48020 23719
rect 47980 23633 48020 23668
rect 47979 23624 48021 23633
rect 47979 23584 47980 23624
rect 48020 23584 48021 23624
rect 47979 23575 48021 23584
rect 47692 23071 47732 23080
rect 48556 23060 48596 24247
rect 48843 24044 48885 24053
rect 48843 24004 48844 24044
rect 48884 24004 48885 24044
rect 48843 23995 48885 24004
rect 48651 23288 48693 23297
rect 48651 23248 48652 23288
rect 48692 23248 48693 23288
rect 48651 23239 48693 23248
rect 48844 23288 48884 23995
rect 48844 23239 48884 23248
rect 47020 23020 47156 23060
rect 48460 23020 48596 23060
rect 46636 20719 46676 20728
rect 46731 20768 46773 20777
rect 46731 20728 46732 20768
rect 46772 20728 46773 20768
rect 46731 20719 46773 20728
rect 46348 20634 46388 20719
rect 44372 20560 44660 20600
rect 44332 20551 44372 20560
rect 44332 20012 44372 20021
rect 44236 19972 44332 20012
rect 44332 19963 44372 19972
rect 44523 20012 44565 20021
rect 44523 19972 44524 20012
rect 44564 19972 44565 20012
rect 44523 19963 44565 19972
rect 44139 19928 44181 19937
rect 44139 19888 44140 19928
rect 44180 19888 44181 19928
rect 44139 19879 44181 19888
rect 44524 19928 44564 19963
rect 43851 19844 43893 19853
rect 43851 19804 43852 19844
rect 43892 19804 43893 19844
rect 43851 19795 43893 19804
rect 43852 19710 43892 19795
rect 44140 19256 44180 19879
rect 44524 19877 44564 19888
rect 44620 19676 44660 20560
rect 45620 20560 45908 20600
rect 45580 20551 45620 20560
rect 44811 20264 44853 20273
rect 44811 20224 44812 20264
rect 44852 20224 44853 20264
rect 44811 20215 44853 20224
rect 44715 19928 44757 19937
rect 44715 19888 44716 19928
rect 44756 19888 44757 19928
rect 44715 19879 44757 19888
rect 44716 19794 44756 19879
rect 44620 19636 44756 19676
rect 44140 19207 44180 19216
rect 44331 19256 44373 19265
rect 44331 19216 44332 19256
rect 44372 19216 44373 19256
rect 44331 19207 44373 19216
rect 43756 19172 43796 19181
rect 43796 19132 44084 19172
rect 43756 19123 43796 19132
rect 43660 18964 43892 19004
rect 43564 18535 43604 18544
rect 43659 18584 43701 18593
rect 43659 18544 43660 18584
rect 43700 18544 43701 18584
rect 43659 18535 43701 18544
rect 43756 18584 43796 18595
rect 43660 18450 43700 18535
rect 43756 18509 43796 18544
rect 43755 18500 43797 18509
rect 43755 18460 43756 18500
rect 43796 18460 43797 18500
rect 43755 18451 43797 18460
rect 43564 17744 43604 17753
rect 43564 16904 43604 17704
rect 43660 16904 43700 16913
rect 43564 16864 43660 16904
rect 43660 16855 43700 16864
rect 43852 16745 43892 18964
rect 44044 18752 44084 19132
rect 44044 18703 44084 18712
rect 43947 18668 43989 18677
rect 43947 18628 43948 18668
rect 43988 18628 43989 18668
rect 43947 18619 43989 18628
rect 43948 18584 43988 18619
rect 43948 17837 43988 18544
rect 44043 18584 44085 18593
rect 44140 18584 44180 18593
rect 44043 18544 44044 18584
rect 44084 18544 44140 18584
rect 44043 18535 44085 18544
rect 44140 18535 44180 18544
rect 44235 18584 44277 18593
rect 44235 18544 44236 18584
rect 44276 18544 44277 18584
rect 44235 18535 44277 18544
rect 44236 18450 44276 18535
rect 44235 18332 44277 18341
rect 44235 18292 44236 18332
rect 44276 18292 44277 18332
rect 44235 18283 44277 18292
rect 43947 17828 43989 17837
rect 43947 17788 43948 17828
rect 43988 17788 43989 17828
rect 43947 17779 43989 17788
rect 44139 17744 44181 17753
rect 44139 17704 44140 17744
rect 44180 17704 44181 17744
rect 44139 17695 44181 17704
rect 44140 17156 44180 17695
rect 44140 17107 44180 17116
rect 44044 17072 44084 17081
rect 44044 16913 44084 17032
rect 44236 17072 44276 18283
rect 44332 17744 44372 19207
rect 44619 18920 44661 18929
rect 44619 18880 44620 18920
rect 44660 18880 44661 18920
rect 44619 18871 44661 18880
rect 44428 18584 44468 18593
rect 44428 18425 44468 18544
rect 44523 18584 44565 18593
rect 44523 18544 44524 18584
rect 44564 18544 44565 18584
rect 44523 18535 44565 18544
rect 44620 18584 44660 18871
rect 44524 18450 44564 18535
rect 44620 18425 44660 18544
rect 44427 18416 44469 18425
rect 44427 18376 44428 18416
rect 44468 18376 44469 18416
rect 44427 18367 44469 18376
rect 44619 18416 44661 18425
rect 44619 18376 44620 18416
rect 44660 18376 44661 18416
rect 44619 18367 44661 18376
rect 44716 18089 44756 19636
rect 44715 18080 44757 18089
rect 44715 18040 44716 18080
rect 44756 18040 44757 18080
rect 44715 18031 44757 18040
rect 44428 17744 44468 17753
rect 44332 17704 44428 17744
rect 44428 17695 44468 17704
rect 44043 16904 44085 16913
rect 44043 16864 44044 16904
rect 44084 16864 44085 16904
rect 44043 16855 44085 16864
rect 43851 16736 43893 16745
rect 43851 16696 43852 16736
rect 43892 16696 43893 16736
rect 43851 16687 43893 16696
rect 43660 16232 43700 16241
rect 43700 16192 43796 16232
rect 43660 16183 43700 16192
rect 43659 15392 43701 15401
rect 43659 15352 43660 15392
rect 43700 15352 43701 15392
rect 43659 15343 43701 15352
rect 43756 15392 43796 16192
rect 44236 15401 44276 17032
rect 44524 16988 44564 16997
rect 44524 16745 44564 16948
rect 44715 16904 44757 16913
rect 44715 16864 44716 16904
rect 44756 16864 44757 16904
rect 44715 16855 44757 16864
rect 44716 16770 44756 16855
rect 44523 16736 44565 16745
rect 44523 16696 44524 16736
rect 44564 16696 44565 16736
rect 44523 16687 44565 16696
rect 44524 16232 44564 16241
rect 44524 16073 44564 16192
rect 44331 16064 44373 16073
rect 44331 16024 44332 16064
rect 44372 16024 44373 16064
rect 44331 16015 44373 16024
rect 44523 16064 44565 16073
rect 44523 16024 44524 16064
rect 44564 16024 44565 16064
rect 44523 16015 44565 16024
rect 43756 15343 43796 15352
rect 44235 15392 44277 15401
rect 44235 15352 44236 15392
rect 44276 15352 44277 15392
rect 44235 15343 44277 15352
rect 43468 15184 43604 15224
rect 42700 14848 43028 14888
rect 43084 14848 43316 14888
rect 42603 14720 42645 14729
rect 42603 14680 42604 14720
rect 42644 14680 42645 14720
rect 42603 14671 42645 14680
rect 42603 14216 42645 14225
rect 42603 14176 42604 14216
rect 42644 14176 42645 14216
rect 42603 14167 42645 14176
rect 42604 13796 42644 14167
rect 42700 13964 42740 14848
rect 42795 14720 42837 14729
rect 42795 14680 42796 14720
rect 42836 14680 42837 14720
rect 42795 14671 42837 14680
rect 42988 14720 43028 14848
rect 42988 14671 43028 14680
rect 43083 14720 43125 14729
rect 43083 14680 43084 14720
rect 43124 14680 43125 14720
rect 43083 14671 43125 14680
rect 43276 14720 43316 14848
rect 43276 14671 43316 14680
rect 43371 14720 43413 14729
rect 43371 14680 43372 14720
rect 43412 14680 43413 14720
rect 43371 14671 43413 14680
rect 43468 14720 43508 14729
rect 42796 14586 42836 14671
rect 43084 14586 43124 14671
rect 43372 14586 43412 14671
rect 42892 14552 42932 14561
rect 42932 14512 43028 14552
rect 42892 14503 42932 14512
rect 42700 13924 42836 13964
rect 42700 13796 42740 13805
rect 42604 13756 42700 13796
rect 42700 13747 42740 13756
rect 42796 13460 42836 13924
rect 42603 13376 42645 13385
rect 42603 13336 42604 13376
rect 42644 13336 42645 13376
rect 42603 13327 42645 13336
rect 42412 12940 42548 12980
rect 42315 12872 42357 12881
rect 42315 12832 42316 12872
rect 42356 12832 42357 12872
rect 42315 12823 42357 12832
rect 42220 12487 42260 12496
rect 42411 12536 42453 12545
rect 42411 12496 42412 12536
rect 42452 12496 42453 12536
rect 42411 12487 42453 12496
rect 42315 12284 42357 12293
rect 42315 12244 42316 12284
rect 42356 12244 42357 12284
rect 42315 12235 42357 12244
rect 42316 12150 42356 12235
rect 42412 12041 42452 12487
rect 42411 12032 42453 12041
rect 42411 11992 42412 12032
rect 42452 11992 42453 12032
rect 42411 11983 42453 11992
rect 42124 11864 42164 11873
rect 42164 11824 42356 11864
rect 42124 11815 42164 11824
rect 42124 11696 42164 11705
rect 42028 11656 42124 11696
rect 41932 11192 41972 11656
rect 42124 11369 42164 11656
rect 42316 11696 42356 11824
rect 42316 11647 42356 11656
rect 42123 11360 42165 11369
rect 42123 11320 42124 11360
rect 42164 11320 42165 11360
rect 42123 11311 42165 11320
rect 42508 11201 42548 12940
rect 42123 11192 42165 11201
rect 41932 11152 42068 11192
rect 41836 11024 41876 11033
rect 41740 10984 41836 11024
rect 41548 10865 41588 10984
rect 41836 10975 41876 10984
rect 41932 11024 41972 11033
rect 41547 10856 41589 10865
rect 41547 10816 41548 10856
rect 41588 10816 41589 10856
rect 41547 10807 41589 10816
rect 41740 10436 41780 10445
rect 41932 10436 41972 10984
rect 42028 10781 42068 11152
rect 42123 11152 42124 11192
rect 42164 11152 42165 11192
rect 42123 11143 42165 11152
rect 42507 11192 42549 11201
rect 42507 11152 42508 11192
rect 42548 11152 42549 11192
rect 42507 11143 42549 11152
rect 42027 10772 42069 10781
rect 42027 10732 42028 10772
rect 42068 10732 42069 10772
rect 42027 10723 42069 10732
rect 42124 10445 42164 11143
rect 42412 11024 42452 11033
rect 42220 10856 42260 10865
rect 42412 10856 42452 10984
rect 42604 11024 42644 13327
rect 42796 13217 42836 13420
rect 42892 13796 42932 13805
rect 42700 13208 42740 13217
rect 42700 13049 42740 13168
rect 42795 13208 42837 13217
rect 42795 13168 42796 13208
rect 42836 13168 42837 13208
rect 42795 13159 42837 13168
rect 42892 13208 42932 13756
rect 42988 13208 43028 14512
rect 43468 14468 43508 14680
rect 43276 14428 43508 14468
rect 43179 14132 43221 14141
rect 43179 14092 43180 14132
rect 43220 14092 43221 14132
rect 43179 14083 43221 14092
rect 43180 13998 43220 14083
rect 43276 14048 43316 14428
rect 43564 14141 43604 15184
rect 43371 14132 43413 14141
rect 43371 14092 43372 14132
rect 43412 14092 43413 14132
rect 43371 14083 43413 14092
rect 43563 14132 43605 14141
rect 43563 14092 43564 14132
rect 43604 14092 43605 14132
rect 43563 14083 43605 14092
rect 43276 13469 43316 14008
rect 43275 13460 43317 13469
rect 43275 13420 43276 13460
rect 43316 13420 43317 13460
rect 43275 13411 43317 13420
rect 43084 13208 43124 13217
rect 42988 13168 43084 13208
rect 42892 13159 42932 13168
rect 43084 13159 43124 13168
rect 42699 13040 42741 13049
rect 42699 13000 42700 13040
rect 42740 13000 42741 13040
rect 42699 12991 42741 13000
rect 42987 12872 43029 12881
rect 43372 12872 43412 14083
rect 43564 14048 43604 14083
rect 43564 13998 43604 14008
rect 43467 13712 43509 13721
rect 43467 13672 43468 13712
rect 43508 13672 43509 13712
rect 43467 13663 43509 13672
rect 43468 13208 43508 13663
rect 43468 13159 43508 13168
rect 43660 13049 43700 15343
rect 44332 14141 44372 16015
rect 44331 14132 44373 14141
rect 44331 14092 44332 14132
rect 44372 14092 44373 14132
rect 44331 14083 44373 14092
rect 43852 13880 43892 13889
rect 43852 13721 43892 13840
rect 43851 13712 43893 13721
rect 43851 13672 43852 13712
rect 43892 13672 43893 13712
rect 43851 13663 43893 13672
rect 44332 13208 44372 14083
rect 43659 13040 43701 13049
rect 43659 13000 43660 13040
rect 43700 13000 43701 13040
rect 43659 12991 43701 13000
rect 42987 12832 42988 12872
rect 43028 12832 43029 12872
rect 42987 12823 43029 12832
rect 43084 12832 43412 12872
rect 42796 12368 42836 12377
rect 42700 12328 42796 12368
rect 42700 11696 42740 12328
rect 42796 12319 42836 12328
rect 42700 11647 42740 11656
rect 42604 10975 42644 10984
rect 42260 10816 42452 10856
rect 42220 10807 42260 10816
rect 42507 10772 42549 10781
rect 42507 10732 42508 10772
rect 42548 10732 42549 10772
rect 42507 10723 42549 10732
rect 42508 10638 42548 10723
rect 41780 10396 41972 10436
rect 42123 10436 42165 10445
rect 42123 10396 42124 10436
rect 42164 10396 42165 10436
rect 41740 10109 41780 10396
rect 42123 10387 42165 10396
rect 42124 10268 42164 10387
rect 42124 10219 42164 10228
rect 41739 10100 41781 10109
rect 41653 10060 41740 10100
rect 41780 10060 41781 10100
rect 41653 9932 41693 10060
rect 41739 10051 41781 10060
rect 42219 10100 42261 10109
rect 42219 10060 42220 10100
rect 42260 10060 42261 10100
rect 42219 10051 42261 10060
rect 41835 10016 41877 10025
rect 41835 9976 41836 10016
rect 41876 9976 41877 10016
rect 41835 9967 41877 9976
rect 41644 9892 41693 9932
rect 41355 9596 41397 9605
rect 41355 9556 41356 9596
rect 41396 9556 41397 9596
rect 41355 9547 41397 9556
rect 40876 9463 40916 9472
rect 41644 9512 41684 9892
rect 41739 9848 41781 9857
rect 41739 9808 41740 9848
rect 41780 9808 41781 9848
rect 41739 9799 41781 9808
rect 41644 9463 41684 9472
rect 41740 9512 41780 9799
rect 41740 9463 41780 9472
rect 39476 9304 39956 9344
rect 41452 9344 41492 9353
rect 39436 9295 39476 9304
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 41452 8681 41492 9304
rect 41547 9260 41589 9269
rect 41547 9220 41548 9260
rect 41588 9220 41589 9260
rect 41547 9211 41589 9220
rect 41451 8672 41493 8681
rect 41451 8632 41452 8672
rect 41492 8632 41493 8672
rect 41451 8623 41493 8632
rect 41548 8588 41588 9211
rect 41836 8765 41876 9967
rect 41931 9596 41973 9605
rect 41931 9556 41932 9596
rect 41972 9556 41973 9596
rect 41931 9547 41973 9556
rect 41932 9512 41972 9547
rect 41932 9461 41972 9472
rect 42124 9512 42164 9521
rect 41932 9344 41972 9353
rect 42124 9344 42164 9472
rect 42220 9512 42260 10051
rect 42316 10016 42356 10027
rect 42316 9941 42356 9976
rect 42315 9932 42357 9941
rect 42315 9892 42316 9932
rect 42356 9892 42357 9932
rect 42315 9883 42357 9892
rect 42795 9680 42837 9689
rect 42795 9640 42796 9680
rect 42836 9640 42837 9680
rect 42795 9631 42837 9640
rect 42220 9463 42260 9472
rect 42412 9512 42452 9521
rect 42604 9512 42644 9521
rect 42452 9472 42604 9512
rect 42412 9463 42452 9472
rect 42604 9463 42644 9472
rect 42699 9512 42741 9521
rect 42699 9472 42700 9512
rect 42740 9472 42741 9512
rect 42699 9463 42741 9472
rect 42796 9512 42836 9631
rect 42988 9605 43028 12823
rect 43084 10865 43124 12832
rect 44332 11705 44372 13168
rect 44620 14048 44660 14057
rect 44427 13040 44469 13049
rect 44427 13000 44428 13040
rect 44468 13000 44469 13040
rect 44427 12991 44469 13000
rect 43563 11696 43605 11705
rect 43563 11656 43564 11696
rect 43604 11656 43605 11696
rect 43563 11647 43605 11656
rect 44331 11696 44373 11705
rect 44331 11656 44332 11696
rect 44372 11656 44373 11696
rect 44331 11647 44373 11656
rect 43564 11562 43604 11647
rect 43947 11276 43989 11285
rect 43947 11236 43948 11276
rect 43988 11236 43989 11276
rect 43947 11227 43989 11236
rect 43467 11192 43509 11201
rect 43467 11152 43468 11192
rect 43508 11152 43509 11192
rect 43467 11143 43509 11152
rect 43851 11192 43893 11201
rect 43851 11152 43852 11192
rect 43892 11152 43893 11192
rect 43851 11143 43893 11152
rect 43276 11024 43316 11033
rect 43083 10856 43125 10865
rect 43083 10816 43084 10856
rect 43124 10816 43125 10856
rect 43083 10807 43125 10816
rect 43084 10193 43124 10807
rect 43083 10184 43125 10193
rect 43083 10144 43084 10184
rect 43124 10144 43125 10184
rect 43083 10135 43125 10144
rect 43276 9941 43316 10984
rect 43468 11024 43508 11143
rect 43468 10975 43508 10984
rect 43660 11024 43700 11033
rect 43372 10856 43412 10865
rect 43660 10856 43700 10984
rect 43412 10816 43700 10856
rect 43756 11024 43796 11033
rect 43372 10807 43412 10816
rect 43756 10436 43796 10984
rect 43660 10396 43796 10436
rect 43467 10184 43509 10193
rect 43467 10144 43468 10184
rect 43508 10144 43509 10184
rect 43467 10135 43509 10144
rect 43468 10050 43508 10135
rect 43660 10109 43700 10396
rect 43852 10352 43892 11143
rect 43948 11024 43988 11227
rect 43948 10975 43988 10984
rect 44140 11024 44180 11033
rect 43948 10856 43988 10865
rect 44140 10856 44180 10984
rect 43988 10816 44180 10856
rect 43948 10807 43988 10816
rect 43756 10312 43892 10352
rect 44140 10352 44180 10361
rect 44180 10312 44372 10352
rect 43756 10184 43796 10312
rect 44140 10303 44180 10312
rect 43756 10135 43796 10144
rect 44332 10184 44372 10312
rect 44428 10268 44468 12991
rect 44620 12041 44660 14008
rect 44812 12713 44852 20215
rect 45003 20180 45045 20189
rect 45003 20140 45004 20180
rect 45044 20140 45045 20180
rect 45003 20131 45045 20140
rect 45004 19265 45044 20131
rect 45195 20096 45237 20105
rect 45195 20056 45196 20096
rect 45236 20056 45237 20096
rect 45195 20047 45237 20056
rect 45100 19844 45140 19853
rect 45003 19256 45045 19265
rect 45003 19216 45004 19256
rect 45044 19216 45045 19256
rect 45003 19207 45045 19216
rect 45004 19122 45044 19207
rect 45100 18509 45140 19804
rect 45099 18500 45141 18509
rect 45099 18460 45100 18500
rect 45140 18460 45141 18500
rect 45099 18451 45141 18460
rect 44907 18080 44949 18089
rect 44907 18040 44908 18080
rect 44948 18040 44949 18080
rect 44907 18031 44949 18040
rect 44908 16988 44948 18031
rect 44908 16939 44948 16948
rect 45099 16820 45141 16829
rect 45099 16780 45100 16820
rect 45140 16780 45141 16820
rect 45099 16771 45141 16780
rect 45100 16686 45140 16771
rect 45196 15233 45236 20047
rect 45291 20012 45333 20021
rect 45291 19972 45292 20012
rect 45332 19972 45333 20012
rect 45291 19963 45333 19972
rect 45676 20012 45716 20021
rect 45292 19878 45332 19963
rect 45484 19844 45524 19853
rect 45484 18677 45524 19804
rect 45579 18752 45621 18761
rect 45579 18712 45580 18752
rect 45620 18712 45621 18752
rect 45579 18703 45621 18712
rect 45483 18668 45525 18677
rect 45483 18628 45484 18668
rect 45524 18628 45525 18668
rect 45483 18619 45525 18628
rect 45483 18416 45525 18425
rect 45580 18416 45620 18703
rect 45483 18376 45484 18416
rect 45524 18376 45620 18416
rect 45483 18367 45525 18376
rect 45291 18164 45333 18173
rect 45291 18124 45292 18164
rect 45332 18124 45333 18164
rect 45291 18115 45333 18124
rect 45195 15224 45237 15233
rect 45195 15184 45196 15224
rect 45236 15184 45237 15224
rect 45195 15175 45237 15184
rect 45100 14888 45140 14897
rect 45004 14048 45044 14057
rect 45100 14048 45140 14848
rect 45292 14804 45332 18115
rect 45388 17072 45428 17081
rect 45388 16913 45428 17032
rect 45387 16904 45429 16913
rect 45387 16864 45388 16904
rect 45428 16864 45429 16904
rect 45387 16855 45429 16864
rect 45484 16073 45524 18367
rect 45676 18089 45716 19972
rect 46635 20012 46677 20021
rect 46635 19972 46636 20012
rect 46676 19972 46677 20012
rect 46635 19963 46677 19972
rect 46348 19172 46388 19181
rect 46388 19132 46484 19172
rect 46348 19123 46388 19132
rect 46156 19088 46196 19097
rect 46156 18761 46196 19048
rect 46155 18752 46197 18761
rect 46155 18712 46156 18752
rect 46196 18712 46197 18752
rect 46155 18703 46197 18712
rect 46155 18584 46197 18593
rect 46155 18544 46156 18584
rect 46196 18544 46197 18584
rect 46155 18535 46197 18544
rect 46348 18584 46388 18593
rect 46156 18450 46196 18535
rect 46251 18416 46293 18425
rect 46251 18376 46252 18416
rect 46292 18376 46293 18416
rect 46251 18367 46293 18376
rect 45867 18332 45909 18341
rect 45867 18292 45868 18332
rect 45908 18292 45909 18332
rect 45867 18283 45909 18292
rect 45675 18080 45717 18089
rect 45675 18040 45676 18080
rect 45716 18040 45717 18080
rect 45675 18031 45717 18040
rect 45868 18005 45908 18283
rect 46252 18282 46292 18367
rect 46348 18332 46388 18544
rect 46444 18509 46484 19132
rect 46443 18500 46485 18509
rect 46443 18460 46444 18500
rect 46484 18460 46485 18500
rect 46443 18451 46485 18460
rect 46348 18292 46484 18332
rect 45963 18164 46005 18173
rect 45963 18124 45964 18164
rect 46004 18124 46005 18164
rect 45963 18115 46005 18124
rect 45867 17996 45909 18005
rect 45867 17956 45868 17996
rect 45908 17956 45909 17996
rect 45867 17947 45909 17956
rect 45964 17669 46004 18115
rect 46347 17996 46389 18005
rect 46347 17956 46348 17996
rect 46388 17956 46389 17996
rect 46347 17947 46389 17956
rect 46348 17862 46388 17947
rect 46060 17744 46100 17753
rect 46156 17744 46196 17753
rect 45963 17660 46005 17669
rect 45963 17620 45964 17660
rect 46004 17620 46005 17660
rect 45963 17611 46005 17620
rect 45580 17576 45620 17585
rect 45580 16157 45620 17536
rect 45772 17156 45812 17165
rect 46060 17156 46100 17704
rect 46155 17704 46156 17744
rect 46155 17695 46196 17704
rect 46348 17744 46388 17755
rect 46155 17585 46195 17695
rect 46348 17669 46388 17704
rect 46347 17660 46389 17669
rect 46347 17620 46348 17660
rect 46388 17620 46389 17660
rect 46347 17611 46389 17620
rect 46444 17585 46484 18292
rect 46539 18248 46581 18257
rect 46539 18208 46540 18248
rect 46580 18208 46581 18248
rect 46539 18199 46581 18208
rect 46540 17828 46580 18199
rect 46540 17779 46580 17788
rect 46155 17576 46197 17585
rect 46155 17536 46156 17576
rect 46196 17536 46197 17576
rect 46155 17527 46197 17536
rect 46443 17576 46485 17585
rect 46443 17536 46444 17576
rect 46484 17536 46485 17576
rect 46443 17527 46485 17536
rect 46636 17240 46676 19963
rect 46828 19928 46868 19937
rect 46732 19888 46828 19928
rect 46732 19256 46772 19888
rect 46828 19879 46868 19888
rect 47020 19517 47060 23020
rect 48172 22448 48212 22457
rect 48076 22408 48172 22448
rect 47212 21608 47252 21617
rect 47212 20777 47252 21568
rect 47691 21356 47733 21365
rect 47691 21316 47692 21356
rect 47732 21316 47733 21356
rect 47691 21307 47733 21316
rect 47211 20768 47253 20777
rect 47211 20728 47212 20768
rect 47252 20728 47253 20768
rect 47211 20719 47253 20728
rect 47595 20768 47637 20777
rect 47595 20728 47596 20768
rect 47636 20728 47637 20768
rect 47595 20719 47637 20728
rect 47692 20768 47732 21307
rect 47692 20719 47732 20728
rect 48076 20768 48116 22408
rect 48172 22399 48212 22408
rect 48363 21524 48405 21533
rect 48460 21524 48500 23020
rect 48555 22280 48597 22289
rect 48555 22240 48556 22280
rect 48596 22240 48597 22280
rect 48555 22231 48597 22240
rect 48652 22280 48692 23239
rect 48747 23204 48789 23213
rect 48747 23164 48748 23204
rect 48788 23164 48789 23204
rect 48747 23155 48789 23164
rect 48652 22231 48692 22240
rect 48748 22280 48788 23155
rect 48940 22289 48980 26095
rect 49228 25985 49268 26104
rect 49227 25976 49269 25985
rect 49227 25936 49228 25976
rect 49268 25936 49269 25976
rect 49227 25927 49269 25936
rect 49420 25733 49460 28624
rect 49515 27572 49557 27581
rect 49515 27532 49516 27572
rect 49556 27532 49557 27572
rect 49515 27523 49557 27532
rect 49516 27068 49556 27523
rect 49516 27019 49556 27028
rect 49516 26648 49556 26657
rect 49516 26405 49556 26608
rect 49515 26396 49557 26405
rect 49515 26356 49516 26396
rect 49556 26356 49557 26396
rect 49515 26347 49557 26356
rect 49419 25724 49461 25733
rect 49419 25684 49420 25724
rect 49460 25684 49461 25724
rect 49419 25675 49461 25684
rect 49612 25556 49652 29044
rect 49803 29000 49845 29009
rect 49803 28960 49804 29000
rect 49844 28960 49845 29000
rect 49803 28951 49845 28960
rect 49804 28866 49844 28951
rect 49996 28757 50036 29044
rect 50380 29009 50420 29128
rect 50476 29168 50516 29791
rect 50572 29681 50612 29800
rect 50667 29840 50709 29849
rect 50667 29800 50668 29840
rect 50708 29800 50709 29840
rect 50667 29791 50709 29800
rect 50668 29706 50708 29791
rect 50571 29672 50613 29681
rect 50571 29632 50572 29672
rect 50612 29632 50613 29672
rect 50571 29623 50613 29632
rect 50764 29168 50804 30379
rect 50860 29924 50900 30724
rect 51147 30764 51189 30773
rect 51147 30724 51148 30764
rect 51188 30724 51189 30764
rect 51147 30715 51189 30724
rect 51723 30764 51765 30773
rect 51723 30724 51724 30764
rect 51764 30724 51765 30764
rect 51723 30715 51765 30724
rect 50956 30680 50996 30689
rect 50956 30092 50996 30640
rect 51148 30680 51188 30715
rect 51148 30629 51188 30640
rect 51340 30680 51380 30689
rect 51244 30437 51284 30522
rect 51243 30428 51285 30437
rect 51243 30388 51244 30428
rect 51284 30388 51285 30428
rect 51340 30428 51380 30640
rect 51532 30605 51572 30690
rect 51820 30689 51860 31144
rect 51819 30680 51861 30689
rect 51819 30640 51820 30680
rect 51860 30640 51861 30680
rect 51819 30631 51861 30640
rect 51531 30596 51573 30605
rect 51531 30556 51532 30596
rect 51572 30556 51573 30596
rect 51531 30547 51573 30556
rect 51916 30596 51956 31387
rect 53452 31361 53492 32143
rect 54412 32117 54452 32152
rect 54604 32192 54644 32201
rect 54411 32108 54453 32117
rect 54411 32068 54412 32108
rect 54452 32068 54453 32108
rect 54411 32059 54453 32068
rect 53547 32024 53589 32033
rect 53547 31984 53548 32024
rect 53588 31984 53589 32024
rect 53547 31975 53589 31984
rect 53548 31890 53588 31975
rect 52107 31352 52149 31361
rect 52107 31312 52108 31352
rect 52148 31312 52149 31352
rect 52107 31303 52149 31312
rect 53164 31352 53204 31361
rect 52108 30857 52148 31303
rect 52780 31268 52820 31277
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 52107 30848 52149 30857
rect 52107 30808 52108 30848
rect 52148 30808 52149 30848
rect 52107 30799 52149 30808
rect 52108 30714 52148 30799
rect 52203 30596 52245 30605
rect 51956 30556 52052 30596
rect 51916 30547 51956 30556
rect 51627 30512 51669 30521
rect 51627 30472 51628 30512
rect 51668 30472 51669 30512
rect 51627 30463 51669 30472
rect 51340 30388 51572 30428
rect 51243 30379 51285 30388
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 50956 30043 50996 30052
rect 50860 29884 50996 29924
rect 50860 29168 50900 29177
rect 50764 29128 50860 29168
rect 50476 29119 50516 29128
rect 50860 29119 50900 29128
rect 50956 29168 50996 29884
rect 51244 29756 51284 29765
rect 51052 29336 51092 29345
rect 51244 29336 51284 29716
rect 51532 29681 51572 30388
rect 51628 29840 51668 30463
rect 51724 30437 51764 30522
rect 51723 30428 51765 30437
rect 51723 30388 51724 30428
rect 51764 30388 51765 30428
rect 51723 30379 51765 30388
rect 51723 30260 51765 30269
rect 51723 30220 51724 30260
rect 51764 30220 51765 30260
rect 51723 30211 51765 30220
rect 51628 29791 51668 29800
rect 51531 29672 51573 29681
rect 51531 29632 51532 29672
rect 51572 29632 51573 29672
rect 51531 29623 51573 29632
rect 51092 29296 51284 29336
rect 51052 29287 51092 29296
rect 50956 29119 50996 29128
rect 51148 29168 51188 29177
rect 51724 29168 51764 30211
rect 51188 29128 51764 29168
rect 51148 29119 51188 29128
rect 50379 29000 50421 29009
rect 50379 28960 50380 29000
rect 50420 28960 50421 29000
rect 50379 28951 50421 28960
rect 50188 28916 50228 28925
rect 50228 28876 50324 28916
rect 50188 28867 50228 28876
rect 49995 28748 50037 28757
rect 49995 28708 49996 28748
rect 50036 28708 50037 28748
rect 49995 28699 50037 28708
rect 50187 28496 50229 28505
rect 50187 28456 50188 28496
rect 50228 28456 50229 28496
rect 50187 28447 50229 28456
rect 49995 28328 50037 28337
rect 49995 28288 49996 28328
rect 50036 28288 50037 28328
rect 49995 28279 50037 28288
rect 50188 28328 50228 28447
rect 50188 28279 50228 28288
rect 50284 28328 50324 28876
rect 50955 28832 50997 28841
rect 50955 28792 50956 28832
rect 50996 28792 50997 28832
rect 50955 28783 50997 28792
rect 50956 28412 50996 28783
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 51339 28580 51381 28589
rect 51339 28540 51340 28580
rect 51380 28540 51381 28580
rect 51339 28531 51381 28540
rect 51340 28446 51380 28531
rect 51723 28496 51765 28505
rect 51723 28456 51724 28496
rect 51764 28456 51765 28496
rect 51723 28447 51765 28456
rect 51148 28412 51188 28421
rect 50956 28372 51148 28412
rect 51148 28363 51188 28372
rect 50284 28279 50324 28288
rect 50475 28328 50517 28337
rect 50475 28288 50476 28328
rect 50516 28288 50517 28328
rect 50475 28279 50517 28288
rect 50572 28328 50612 28339
rect 49996 28194 50036 28279
rect 50476 28194 50516 28279
rect 50572 28253 50612 28288
rect 50668 28328 50708 28337
rect 50571 28244 50613 28253
rect 50571 28204 50572 28244
rect 50612 28204 50613 28244
rect 50571 28195 50613 28204
rect 50668 28169 50708 28288
rect 50763 28328 50805 28337
rect 51243 28328 51285 28337
rect 51628 28328 51668 28337
rect 50763 28288 50764 28328
rect 50804 28288 50900 28328
rect 50763 28279 50805 28288
rect 50764 28194 50804 28279
rect 50091 28160 50133 28169
rect 50091 28120 50092 28160
rect 50132 28120 50133 28160
rect 50091 28111 50133 28120
rect 50667 28160 50709 28169
rect 50667 28120 50668 28160
rect 50708 28120 50709 28160
rect 50667 28111 50709 28120
rect 50092 28026 50132 28111
rect 50091 27656 50133 27665
rect 50091 27616 50092 27656
rect 50132 27616 50133 27656
rect 50091 27607 50133 27616
rect 50092 26144 50132 27607
rect 50571 27572 50613 27581
rect 50571 27532 50572 27572
rect 50612 27532 50613 27572
rect 50571 27523 50613 27532
rect 50398 26993 50438 26998
rect 50397 26984 50439 26993
rect 50572 26984 50612 27523
rect 50397 26944 50398 26984
rect 50438 26944 50439 26984
rect 50397 26935 50439 26944
rect 50564 26944 50612 26984
rect 50398 26903 50438 26935
rect 50398 26854 50438 26863
rect 50564 26900 50604 26944
rect 50564 26860 50612 26900
rect 50572 26827 50612 26860
rect 50188 26648 50228 26657
rect 50283 26648 50325 26657
rect 50228 26608 50284 26648
rect 50324 26608 50325 26648
rect 50188 26599 50228 26608
rect 50283 26599 50325 26608
rect 50092 26095 50132 26104
rect 49995 25724 50037 25733
rect 49995 25684 49996 25724
rect 50036 25684 50037 25724
rect 49995 25675 50037 25684
rect 49420 25516 49652 25556
rect 49227 23960 49269 23969
rect 49227 23920 49228 23960
rect 49268 23920 49269 23960
rect 49227 23911 49269 23920
rect 49228 23792 49268 23911
rect 49228 23743 49268 23752
rect 49420 23060 49460 25516
rect 49516 25136 49556 25147
rect 49516 25061 49556 25096
rect 49515 25052 49557 25061
rect 49515 25012 49516 25052
rect 49556 25012 49557 25052
rect 49515 25003 49557 25012
rect 49515 24716 49557 24725
rect 49515 24676 49516 24716
rect 49556 24676 49557 24716
rect 49515 24667 49557 24676
rect 49516 23288 49556 24667
rect 49996 24548 50036 25675
rect 50187 25304 50229 25313
rect 50187 25264 50188 25304
rect 50228 25264 50229 25304
rect 50187 25255 50229 25264
rect 50188 24800 50228 25255
rect 50188 24751 50228 24760
rect 49996 24499 50036 24508
rect 50284 24548 50324 26599
rect 50572 25808 50612 26787
rect 50764 26816 50804 26825
rect 50764 26657 50804 26776
rect 50860 26816 50900 28288
rect 51243 28288 51244 28328
rect 51284 28288 51285 28328
rect 51243 28279 51285 28288
rect 51436 28288 51628 28328
rect 50955 28244 50997 28253
rect 50955 28204 50956 28244
rect 50996 28204 50997 28244
rect 50955 28195 50997 28204
rect 50860 26767 50900 26776
rect 50668 26648 50708 26657
rect 50668 26153 50708 26608
rect 50763 26648 50805 26657
rect 50763 26608 50764 26648
rect 50804 26608 50805 26648
rect 50763 26599 50805 26608
rect 50956 26228 50996 28195
rect 51244 27824 51284 28279
rect 51244 27775 51284 27784
rect 51436 27488 51476 28288
rect 51628 28279 51668 28288
rect 51531 27992 51573 28001
rect 51531 27952 51532 27992
rect 51572 27952 51573 27992
rect 51531 27943 51573 27952
rect 51532 27656 51572 27943
rect 51627 27740 51669 27749
rect 51627 27700 51628 27740
rect 51668 27700 51669 27740
rect 51627 27691 51669 27700
rect 51532 27607 51572 27616
rect 51628 27606 51668 27691
rect 51724 27656 51764 28447
rect 51820 28328 51860 28337
rect 51860 28288 51956 28328
rect 51820 28279 51860 28288
rect 51724 27607 51764 27616
rect 51820 27656 51860 27665
rect 51436 27448 51668 27488
rect 51244 27404 51284 27413
rect 51284 27364 51572 27404
rect 51244 27355 51284 27364
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 51148 26816 51188 26825
rect 51148 26321 51188 26776
rect 51436 26816 51476 26825
rect 51436 26657 51476 26776
rect 51532 26816 51572 27364
rect 51532 26767 51572 26776
rect 51435 26648 51477 26657
rect 51435 26608 51436 26648
rect 51476 26608 51477 26648
rect 51435 26599 51477 26608
rect 51147 26312 51189 26321
rect 51147 26272 51148 26312
rect 51188 26272 51189 26312
rect 51628 26312 51668 27448
rect 51820 27245 51860 27616
rect 51819 27236 51861 27245
rect 51819 27196 51820 27236
rect 51860 27196 51861 27236
rect 51819 27187 51861 27196
rect 51820 27068 51860 27077
rect 51916 27068 51956 28288
rect 52012 28169 52052 30556
rect 52203 30556 52204 30596
rect 52244 30556 52245 30596
rect 52203 30547 52245 30556
rect 52108 30428 52148 30437
rect 52108 30269 52148 30388
rect 52107 30260 52149 30269
rect 52107 30220 52108 30260
rect 52148 30220 52149 30260
rect 52107 30211 52149 30220
rect 52204 30092 52244 30547
rect 52780 30521 52820 31228
rect 53164 30932 53204 31312
rect 53451 31352 53493 31361
rect 53451 31312 53452 31352
rect 53492 31312 53493 31352
rect 53451 31303 53493 31312
rect 54027 31352 54069 31361
rect 54027 31312 54028 31352
rect 54068 31312 54069 31352
rect 54027 31303 54069 31312
rect 54028 31218 54068 31303
rect 53164 30892 53300 30932
rect 53260 30554 53300 30892
rect 54508 30680 54548 30689
rect 54604 30680 54644 32152
rect 54700 32192 54740 32320
rect 54700 30848 54740 32152
rect 54796 32192 54836 32201
rect 54796 31949 54836 32152
rect 54892 32192 54932 32203
rect 54892 32117 54932 32152
rect 54891 32108 54933 32117
rect 54891 32068 54892 32108
rect 54932 32068 54933 32108
rect 54891 32059 54933 32068
rect 54795 31940 54837 31949
rect 54795 31900 54796 31940
rect 54836 31900 54837 31940
rect 54795 31891 54837 31900
rect 54700 30808 54932 30848
rect 54548 30640 54644 30680
rect 54699 30680 54741 30689
rect 54699 30640 54700 30680
rect 54740 30640 54741 30680
rect 54508 30631 54548 30640
rect 54699 30631 54741 30640
rect 54796 30680 54836 30689
rect 52299 30512 52341 30521
rect 52299 30472 52300 30512
rect 52340 30472 52341 30512
rect 52299 30463 52341 30472
rect 52779 30512 52821 30521
rect 52779 30472 52780 30512
rect 52820 30472 52821 30512
rect 54700 30546 54740 30631
rect 53260 30505 53300 30514
rect 54507 30512 54549 30521
rect 52779 30463 52821 30472
rect 54507 30472 54508 30512
rect 54548 30472 54549 30512
rect 54507 30463 54549 30472
rect 52300 30378 52340 30463
rect 54508 30378 54548 30463
rect 52491 30176 52533 30185
rect 52491 30136 52492 30176
rect 52532 30136 52533 30176
rect 52491 30127 52533 30136
rect 52108 30052 52244 30092
rect 52011 28160 52053 28169
rect 52011 28120 52012 28160
rect 52052 28120 52053 28160
rect 52011 28111 52053 28120
rect 52012 28001 52052 28111
rect 52011 27992 52053 28001
rect 52011 27952 52012 27992
rect 52052 27952 52053 27992
rect 52011 27943 52053 27952
rect 52011 27740 52053 27749
rect 52011 27700 52012 27740
rect 52052 27700 52053 27740
rect 52011 27691 52053 27700
rect 52012 27606 52052 27691
rect 52108 27488 52148 30052
rect 52492 29849 52532 30127
rect 54796 30092 54836 30640
rect 54796 30043 54836 30052
rect 54795 29924 54837 29933
rect 54795 29884 54796 29924
rect 54836 29884 54837 29924
rect 54795 29875 54837 29884
rect 52491 29840 52533 29849
rect 52491 29800 52492 29840
rect 52532 29800 52533 29840
rect 52491 29791 52533 29800
rect 54123 29840 54165 29849
rect 54123 29800 54124 29840
rect 54164 29800 54165 29840
rect 54123 29791 54165 29800
rect 54796 29840 54836 29875
rect 52492 29706 52532 29791
rect 53643 29672 53685 29681
rect 53643 29632 53644 29672
rect 53684 29632 53685 29672
rect 53643 29623 53685 29632
rect 53644 29538 53684 29623
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 52876 29168 52916 29177
rect 52299 29084 52341 29093
rect 52299 29044 52300 29084
rect 52340 29044 52341 29084
rect 52299 29035 52341 29044
rect 52300 28496 52340 29035
rect 52876 28505 52916 29128
rect 53260 29132 53300 29179
rect 54124 29177 54164 29791
rect 54796 29789 54836 29800
rect 54315 29672 54357 29681
rect 54315 29632 54316 29672
rect 54356 29632 54357 29672
rect 54315 29623 54357 29632
rect 53259 29092 53260 29093
rect 54123 29168 54165 29177
rect 54123 29128 54124 29168
rect 54164 29128 54165 29168
rect 54123 29119 54165 29128
rect 53300 29092 53301 29093
rect 53259 29084 53301 29092
rect 53259 29044 53260 29084
rect 53300 29044 53301 29084
rect 53259 29035 53301 29044
rect 54124 29034 54164 29119
rect 52300 28447 52340 28456
rect 52492 28496 52532 28505
rect 52492 28160 52532 28456
rect 52875 28496 52917 28505
rect 52875 28456 52876 28496
rect 52916 28456 52917 28496
rect 52875 28447 52917 28456
rect 52204 28120 52532 28160
rect 52972 28328 53012 28337
rect 52204 27656 52244 28120
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 52396 27656 52436 27665
rect 52204 27616 52396 27656
rect 52396 27607 52436 27616
rect 51860 27028 51956 27068
rect 52012 27448 52148 27488
rect 51820 27019 51860 27028
rect 52012 26984 52052 27448
rect 52107 27236 52149 27245
rect 52107 27196 52108 27236
rect 52148 27196 52149 27236
rect 52107 27187 52149 27196
rect 52108 27068 52148 27187
rect 52108 27019 52148 27028
rect 51916 26944 52052 26984
rect 51628 26272 51860 26312
rect 51147 26263 51189 26272
rect 50764 26188 50996 26228
rect 51531 26228 51573 26237
rect 51531 26188 51532 26228
rect 51572 26188 51573 26228
rect 50667 26144 50709 26153
rect 50667 26104 50668 26144
rect 50708 26104 50709 26144
rect 50667 26095 50709 26104
rect 50476 25768 50612 25808
rect 50476 24725 50516 25768
rect 50571 25472 50613 25481
rect 50571 25432 50572 25472
rect 50612 25432 50613 25472
rect 50571 25423 50613 25432
rect 50572 25304 50612 25423
rect 50668 25313 50708 25398
rect 50572 25136 50612 25264
rect 50667 25304 50709 25313
rect 50667 25264 50668 25304
rect 50708 25264 50709 25304
rect 50667 25255 50709 25264
rect 50764 25304 50804 26188
rect 51531 26179 51573 26188
rect 51436 26144 51476 26153
rect 50572 25096 50708 25136
rect 50475 24716 50517 24725
rect 50380 24674 50420 24683
rect 50475 24676 50476 24716
rect 50516 24676 50517 24716
rect 50475 24674 50517 24676
rect 50420 24667 50517 24674
rect 50420 24634 50516 24667
rect 50380 24625 50420 24634
rect 50572 24632 50612 24641
rect 50572 24548 50612 24592
rect 50668 24632 50708 25096
rect 50668 24583 50708 24592
rect 50284 24508 50612 24548
rect 50188 24389 50228 24474
rect 49803 24380 49845 24389
rect 49803 24340 49804 24380
rect 49844 24340 49845 24380
rect 49803 24331 49845 24340
rect 50187 24380 50229 24389
rect 50187 24340 50188 24380
rect 50228 24340 50229 24380
rect 50187 24331 50229 24340
rect 49804 23297 49844 24331
rect 50284 24212 50324 24508
rect 50379 24380 50421 24389
rect 50379 24340 50380 24380
rect 50420 24340 50421 24380
rect 50379 24331 50421 24340
rect 50380 24246 50420 24331
rect 50188 24172 50324 24212
rect 49899 23960 49941 23969
rect 49899 23920 49900 23960
rect 49940 23920 49941 23960
rect 49899 23911 49941 23920
rect 49516 23239 49556 23248
rect 49803 23288 49845 23297
rect 49803 23248 49804 23288
rect 49844 23248 49845 23288
rect 49803 23239 49845 23248
rect 49708 23129 49748 23214
rect 49707 23120 49749 23129
rect 49707 23080 49708 23120
rect 49748 23080 49749 23120
rect 49707 23071 49749 23080
rect 49804 23120 49844 23239
rect 49900 23213 49940 23911
rect 49995 23792 50037 23801
rect 49995 23752 49996 23792
rect 50036 23752 50037 23792
rect 49995 23743 50037 23752
rect 49996 23288 50036 23743
rect 49996 23239 50036 23248
rect 49899 23204 49941 23213
rect 49899 23164 49900 23204
rect 49940 23164 49941 23204
rect 49899 23155 49941 23164
rect 49804 23071 49844 23080
rect 49900 23120 49940 23155
rect 49324 23036 49460 23060
rect 49364 23020 49460 23036
rect 49324 22987 49364 22996
rect 49516 22868 49556 22877
rect 49035 22364 49077 22373
rect 49035 22324 49036 22364
rect 49076 22324 49077 22364
rect 49035 22315 49077 22324
rect 48748 22231 48788 22240
rect 48939 22280 48981 22289
rect 48939 22240 48940 22280
rect 48980 22240 48981 22280
rect 48939 22231 48981 22240
rect 48363 21484 48364 21524
rect 48404 21484 48500 21524
rect 48363 21475 48405 21484
rect 48364 21390 48404 21475
rect 48556 21029 48596 22231
rect 49036 22230 49076 22315
rect 49420 22280 49460 22289
rect 49516 22280 49556 22828
rect 49460 22240 49556 22280
rect 49612 22280 49652 22289
rect 49420 22231 49460 22240
rect 48844 22112 48884 22121
rect 48844 21608 48884 22072
rect 49227 22112 49269 22121
rect 49516 22112 49556 22121
rect 49227 22072 49228 22112
rect 49268 22072 49269 22112
rect 49227 22063 49269 22072
rect 49324 22072 49516 22112
rect 49612 22112 49652 22240
rect 49708 22280 49748 23071
rect 49900 23070 49940 23080
rect 50188 23045 50228 24172
rect 50764 23969 50804 25264
rect 50860 26104 51436 26144
rect 50860 25304 50900 26104
rect 51436 26095 51476 26104
rect 51532 26094 51572 26179
rect 51628 26144 51668 26153
rect 50955 25976 50997 25985
rect 50955 25936 50956 25976
rect 50996 25936 50997 25976
rect 50955 25927 50997 25936
rect 50956 25304 50996 25927
rect 51244 25901 51284 25986
rect 51243 25892 51285 25901
rect 51243 25852 51244 25892
rect 51284 25852 51285 25892
rect 51243 25843 51285 25852
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 51436 25472 51476 25481
rect 51052 25304 51092 25313
rect 50956 25264 51052 25304
rect 50860 25255 50900 25264
rect 50955 24884 50997 24893
rect 50955 24844 50956 24884
rect 50996 24844 50997 24884
rect 50955 24835 50997 24844
rect 50859 24380 50901 24389
rect 50859 24340 50860 24380
rect 50900 24340 50901 24380
rect 50859 24331 50901 24340
rect 50763 23960 50805 23969
rect 50763 23920 50764 23960
rect 50804 23920 50805 23960
rect 50763 23911 50805 23920
rect 50571 23792 50613 23801
rect 50571 23752 50572 23792
rect 50612 23752 50613 23792
rect 50571 23743 50613 23752
rect 50764 23792 50804 23801
rect 50572 23658 50612 23743
rect 50764 23633 50804 23752
rect 50860 23792 50900 24331
rect 50860 23743 50900 23752
rect 50380 23624 50420 23633
rect 50667 23624 50709 23633
rect 50420 23584 50516 23624
rect 50380 23575 50420 23584
rect 50379 23372 50421 23381
rect 50379 23332 50380 23372
rect 50420 23332 50421 23372
rect 50379 23323 50421 23332
rect 50284 23120 50324 23148
rect 50380 23120 50420 23323
rect 50476 23213 50516 23584
rect 50667 23584 50668 23624
rect 50708 23584 50709 23624
rect 50764 23624 50810 23633
rect 50956 23624 50996 24835
rect 51052 24464 51092 25264
rect 51244 25304 51284 25313
rect 51436 25304 51476 25432
rect 51284 25264 51476 25304
rect 51244 25255 51284 25264
rect 51148 25220 51188 25229
rect 51148 24641 51188 25180
rect 51339 25136 51381 25145
rect 51339 25096 51340 25136
rect 51380 25096 51381 25136
rect 51339 25087 51381 25096
rect 51147 24632 51189 24641
rect 51147 24592 51148 24632
rect 51188 24592 51189 24632
rect 51147 24583 51189 24592
rect 51340 24548 51380 25087
rect 51628 24641 51668 26104
rect 51723 26144 51765 26153
rect 51723 26104 51724 26144
rect 51764 26104 51765 26144
rect 51723 26095 51765 26104
rect 51724 26010 51764 26095
rect 51820 25985 51860 26272
rect 51916 26060 51956 26944
rect 52972 26825 53012 28288
rect 53163 28160 53205 28169
rect 53163 28120 53164 28160
rect 53204 28120 53205 28160
rect 53163 28111 53205 28120
rect 52012 26816 52052 26825
rect 52012 26573 52052 26776
rect 52204 26816 52244 26825
rect 52204 26657 52244 26776
rect 52971 26816 53013 26825
rect 52971 26776 52972 26816
rect 53012 26776 53013 26816
rect 52971 26767 53013 26776
rect 52203 26648 52245 26657
rect 52203 26608 52204 26648
rect 52244 26608 52245 26648
rect 52203 26599 52245 26608
rect 52011 26564 52053 26573
rect 52011 26524 52012 26564
rect 52052 26524 52053 26564
rect 52011 26515 52053 26524
rect 52012 26237 52052 26515
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 52107 26312 52149 26321
rect 52107 26272 52108 26312
rect 52148 26272 52149 26312
rect 52107 26263 52149 26272
rect 52011 26228 52053 26237
rect 52011 26188 52012 26228
rect 52052 26188 52053 26228
rect 52011 26179 52053 26188
rect 52108 26178 52148 26263
rect 52491 26228 52533 26237
rect 52491 26188 52492 26228
rect 52532 26188 52533 26228
rect 52491 26179 52533 26188
rect 52492 26144 52532 26179
rect 52492 26093 52532 26104
rect 52684 26144 52724 26153
rect 51916 26011 51956 26020
rect 51819 25976 51861 25985
rect 51819 25936 51820 25976
rect 51860 25936 51861 25976
rect 51819 25927 51861 25936
rect 52684 25901 52724 26104
rect 52876 25976 52916 25985
rect 52780 25936 52876 25976
rect 51723 25892 51765 25901
rect 51723 25852 51724 25892
rect 51764 25852 51765 25892
rect 51723 25843 51765 25852
rect 52108 25892 52148 25901
rect 52588 25892 52628 25901
rect 51724 25481 51764 25843
rect 51723 25472 51765 25481
rect 51723 25432 51724 25472
rect 51764 25432 51765 25472
rect 51723 25423 51765 25432
rect 51724 25304 51764 25423
rect 51724 25255 51764 25264
rect 51819 25304 51861 25313
rect 51819 25264 51820 25304
rect 51860 25264 51861 25304
rect 51819 25255 51861 25264
rect 52108 25304 52148 25852
rect 51820 25170 51860 25255
rect 52011 25220 52053 25229
rect 52011 25180 52012 25220
rect 52052 25180 52053 25220
rect 52011 25171 52053 25180
rect 51915 25136 51957 25145
rect 51915 25096 51916 25136
rect 51956 25096 51957 25136
rect 51915 25087 51957 25096
rect 51819 24968 51861 24977
rect 51819 24928 51820 24968
rect 51860 24928 51861 24968
rect 51819 24919 51861 24928
rect 51627 24632 51669 24641
rect 51627 24592 51628 24632
rect 51668 24592 51669 24632
rect 51627 24583 51669 24592
rect 51340 24499 51380 24508
rect 51148 24464 51188 24473
rect 51052 24424 51148 24464
rect 51052 23969 51092 24424
rect 51148 24415 51188 24424
rect 51051 23960 51093 23969
rect 51051 23920 51052 23960
rect 51092 23920 51093 23960
rect 51051 23911 51093 23920
rect 51148 23920 51764 23960
rect 51051 23792 51093 23801
rect 51051 23752 51052 23792
rect 51092 23752 51093 23792
rect 51051 23743 51093 23752
rect 50764 23584 50769 23624
rect 50809 23584 50810 23624
rect 50667 23575 50709 23584
rect 50768 23575 50810 23584
rect 50860 23584 50996 23624
rect 50668 23490 50708 23575
rect 50571 23456 50613 23465
rect 50571 23416 50572 23456
rect 50612 23416 50613 23456
rect 50571 23407 50613 23416
rect 50475 23204 50517 23213
rect 50475 23164 50476 23204
rect 50516 23164 50517 23204
rect 50475 23155 50517 23164
rect 50324 23080 50420 23120
rect 50284 23071 50324 23080
rect 50187 23036 50229 23045
rect 50187 22996 50188 23036
rect 50228 22996 50229 23036
rect 50187 22987 50229 22996
rect 49708 22231 49748 22240
rect 50188 22280 50228 22987
rect 50380 22448 50420 23080
rect 50572 23120 50612 23407
rect 50763 23288 50805 23297
rect 50763 23248 50764 23288
rect 50804 23248 50805 23288
rect 50763 23239 50805 23248
rect 50667 23204 50709 23213
rect 50667 23164 50668 23204
rect 50708 23164 50709 23204
rect 50667 23155 50709 23164
rect 50572 23071 50612 23080
rect 50668 23070 50708 23155
rect 50380 22408 50516 22448
rect 50188 22112 50228 22240
rect 50380 22280 50420 22289
rect 50283 22196 50325 22205
rect 50283 22156 50284 22196
rect 50324 22156 50325 22196
rect 50283 22147 50325 22156
rect 49612 22072 50228 22112
rect 49228 21978 49268 22063
rect 48844 21559 48884 21568
rect 49035 21608 49077 21617
rect 49035 21568 49036 21608
rect 49076 21568 49077 21608
rect 49035 21559 49077 21568
rect 49132 21608 49172 21617
rect 49324 21608 49364 22072
rect 49516 22063 49556 22072
rect 50284 22062 50324 22147
rect 50380 22037 50420 22240
rect 50379 22028 50421 22037
rect 50379 21988 50380 22028
rect 50420 21988 50421 22028
rect 50379 21979 50421 21988
rect 49515 21944 49557 21953
rect 49515 21904 49516 21944
rect 49556 21904 49557 21944
rect 49515 21895 49557 21904
rect 49172 21568 49364 21608
rect 49516 21608 49556 21895
rect 50380 21860 50420 21979
rect 50284 21820 50420 21860
rect 49132 21559 49172 21568
rect 49516 21559 49556 21568
rect 49611 21608 49653 21617
rect 49611 21568 49612 21608
rect 49652 21568 49653 21608
rect 49611 21559 49653 21568
rect 49708 21608 49748 21617
rect 49036 21474 49076 21559
rect 49612 21474 49652 21559
rect 49708 21440 49748 21568
rect 50188 21608 50228 21617
rect 49900 21440 49940 21449
rect 49708 21400 49900 21440
rect 49900 21391 49940 21400
rect 48843 21356 48885 21365
rect 48843 21316 48844 21356
rect 48884 21316 48885 21356
rect 48843 21307 48885 21316
rect 48844 21222 48884 21307
rect 48555 21020 48597 21029
rect 48555 20980 48556 21020
rect 48596 20980 48597 21020
rect 48555 20971 48597 20980
rect 50091 21020 50133 21029
rect 50188 21020 50228 21568
rect 50284 21608 50324 21820
rect 50379 21692 50421 21701
rect 50379 21652 50380 21692
rect 50420 21652 50421 21692
rect 50379 21643 50421 21652
rect 50284 21559 50324 21568
rect 50091 20980 50092 21020
rect 50132 20980 50228 21020
rect 50091 20971 50133 20980
rect 50092 20886 50132 20971
rect 48076 20719 48116 20728
rect 48939 20768 48981 20777
rect 48939 20728 48940 20768
rect 48980 20728 48981 20768
rect 48939 20719 48981 20728
rect 50284 20768 50324 20777
rect 50380 20768 50420 21643
rect 50476 21608 50516 22408
rect 50764 22121 50804 23239
rect 50860 22541 50900 23584
rect 51052 23297 51092 23743
rect 51148 23708 51188 23920
rect 51340 23836 51668 23876
rect 51148 23659 51188 23668
rect 51244 23792 51284 23801
rect 51244 23633 51284 23752
rect 51340 23792 51380 23836
rect 51340 23743 51380 23752
rect 51243 23624 51285 23633
rect 51243 23584 51244 23624
rect 51284 23584 51285 23624
rect 51243 23575 51285 23584
rect 51051 23288 51093 23297
rect 51051 23248 51052 23288
rect 51092 23248 51093 23288
rect 51051 23239 51093 23248
rect 51244 23204 51284 23575
rect 51435 23288 51477 23297
rect 51435 23248 51436 23288
rect 51476 23248 51477 23288
rect 51435 23239 51477 23248
rect 51244 23155 51284 23164
rect 51340 23129 51380 23214
rect 51148 23120 51188 23129
rect 51148 23060 51188 23080
rect 51339 23120 51381 23129
rect 51339 23080 51340 23120
rect 51380 23080 51381 23120
rect 51339 23071 51381 23080
rect 50956 23020 51188 23060
rect 50956 22952 50996 23020
rect 50956 22903 50996 22912
rect 51340 22700 51380 23071
rect 51148 22660 51380 22700
rect 50859 22532 50901 22541
rect 50859 22492 50860 22532
rect 50900 22492 50901 22532
rect 50859 22483 50901 22492
rect 50859 22196 50901 22205
rect 50859 22156 50860 22196
rect 50900 22156 50901 22196
rect 50859 22147 50901 22156
rect 50763 22112 50805 22121
rect 50763 22072 50764 22112
rect 50804 22072 50805 22112
rect 50763 22063 50805 22072
rect 50764 21785 50804 22063
rect 50763 21776 50805 21785
rect 50763 21736 50764 21776
rect 50804 21736 50805 21776
rect 50763 21727 50805 21736
rect 50572 21608 50612 21617
rect 50476 21568 50572 21608
rect 50572 21559 50612 21568
rect 50860 21608 50900 22147
rect 51148 21953 51188 22660
rect 51244 22532 51284 22541
rect 51436 22532 51476 23239
rect 51628 23204 51668 23836
rect 51724 23792 51764 23920
rect 51724 23743 51764 23752
rect 51723 23624 51765 23633
rect 51723 23584 51724 23624
rect 51764 23584 51765 23624
rect 51723 23575 51765 23584
rect 51724 23465 51764 23575
rect 51723 23456 51765 23465
rect 51723 23416 51724 23456
rect 51764 23416 51765 23456
rect 51723 23407 51765 23416
rect 51532 23141 51572 23160
rect 51628 23155 51668 23164
rect 51532 23045 51572 23101
rect 51724 23120 51764 23407
rect 51820 23381 51860 24919
rect 51819 23372 51861 23381
rect 51819 23332 51820 23372
rect 51860 23332 51861 23372
rect 51819 23323 51861 23332
rect 51819 23204 51861 23213
rect 51819 23164 51820 23204
rect 51860 23164 51861 23204
rect 51819 23155 51861 23164
rect 51724 23071 51764 23080
rect 51531 23036 51573 23045
rect 51531 22996 51532 23036
rect 51572 22996 51573 23036
rect 51531 22987 51573 22996
rect 51532 22956 51572 22987
rect 51820 22793 51860 23155
rect 51819 22784 51861 22793
rect 51819 22744 51820 22784
rect 51860 22744 51861 22784
rect 51819 22735 51861 22744
rect 51284 22492 51572 22532
rect 51244 22483 51284 22492
rect 51435 22280 51477 22289
rect 51435 22240 51436 22280
rect 51476 22240 51477 22280
rect 51435 22231 51477 22240
rect 51436 22146 51476 22231
rect 51147 21944 51189 21953
rect 51147 21904 51148 21944
rect 51188 21904 51189 21944
rect 51147 21895 51189 21904
rect 51147 21776 51189 21785
rect 51147 21736 51148 21776
rect 51188 21736 51189 21776
rect 51147 21727 51189 21736
rect 51051 21692 51093 21701
rect 51051 21652 51052 21692
rect 51092 21652 51093 21692
rect 51051 21643 51093 21652
rect 50860 21559 50900 21568
rect 50955 21608 50997 21617
rect 50955 21568 50956 21608
rect 50996 21568 50997 21608
rect 50955 21559 50997 21568
rect 50956 21474 50996 21559
rect 51052 21558 51092 21643
rect 51148 21608 51188 21727
rect 51148 21559 51188 21568
rect 51340 21440 51380 21449
rect 51340 21104 51380 21400
rect 50764 21064 51380 21104
rect 50324 20728 50420 20768
rect 50668 20768 50708 20777
rect 50764 20768 50804 21064
rect 51532 20777 51572 22492
rect 50708 20728 50804 20768
rect 50859 20768 50901 20777
rect 50859 20728 50860 20768
rect 50900 20728 50901 20768
rect 50284 20719 50324 20728
rect 50668 20719 50708 20728
rect 50859 20719 50901 20728
rect 51531 20768 51573 20777
rect 51531 20728 51532 20768
rect 51572 20728 51573 20768
rect 51531 20719 51573 20728
rect 47596 20189 47636 20719
rect 48940 20634 48980 20719
rect 47595 20180 47637 20189
rect 47595 20140 47596 20180
rect 47636 20140 47637 20180
rect 47595 20131 47637 20140
rect 47500 20012 47540 20021
rect 47404 19972 47500 20012
rect 47307 19844 47349 19853
rect 47307 19804 47308 19844
rect 47348 19804 47349 19844
rect 47307 19795 47349 19804
rect 47308 19710 47348 19795
rect 47019 19508 47061 19517
rect 47019 19468 47020 19508
rect 47060 19468 47061 19508
rect 47019 19459 47061 19468
rect 46732 19207 46772 19216
rect 47404 18929 47444 19972
rect 47500 19963 47540 19972
rect 47499 19844 47541 19853
rect 47499 19804 47500 19844
rect 47540 19804 47541 19844
rect 47499 19795 47541 19804
rect 47403 18920 47445 18929
rect 47403 18880 47404 18920
rect 47444 18880 47445 18920
rect 47403 18871 47445 18880
rect 47500 18752 47540 19795
rect 47596 19256 47636 20131
rect 47884 20012 47924 20021
rect 49323 20012 49365 20021
rect 47924 19972 48020 20012
rect 47884 19963 47924 19972
rect 47691 19844 47733 19853
rect 47691 19804 47692 19844
rect 47732 19804 47733 19844
rect 47691 19795 47733 19804
rect 47692 19710 47732 19795
rect 47980 19676 48020 19972
rect 49323 19972 49324 20012
rect 49364 19972 49365 20012
rect 49323 19963 49365 19972
rect 49324 19878 49364 19963
rect 50092 19928 50132 19937
rect 49996 19888 50092 19928
rect 49132 19844 49172 19853
rect 47980 19636 48500 19676
rect 47636 19216 47828 19256
rect 47596 19207 47636 19216
rect 47500 18712 47636 18752
rect 46827 18668 46869 18677
rect 46827 18628 46828 18668
rect 46868 18628 46869 18668
rect 46827 18619 46869 18628
rect 46732 18584 46772 18593
rect 46732 18005 46772 18544
rect 46828 18584 46868 18619
rect 46828 18533 46868 18544
rect 47019 18584 47061 18593
rect 47019 18544 47020 18584
rect 47060 18544 47061 18584
rect 47019 18535 47061 18544
rect 47403 18584 47445 18593
rect 47403 18544 47404 18584
rect 47444 18544 47445 18584
rect 47403 18535 47445 18544
rect 47500 18584 47540 18593
rect 46923 18500 46965 18509
rect 46923 18460 46924 18500
rect 46964 18460 46965 18500
rect 46923 18451 46965 18460
rect 46827 18416 46869 18425
rect 46827 18376 46828 18416
rect 46868 18376 46869 18416
rect 46827 18367 46869 18376
rect 46731 17996 46773 18005
rect 46731 17956 46732 17996
rect 46772 17956 46773 17996
rect 46731 17947 46773 17956
rect 46731 17576 46773 17585
rect 46731 17536 46732 17576
rect 46772 17536 46773 17576
rect 46731 17527 46773 17536
rect 46732 17442 46772 17527
rect 46828 17333 46868 18367
rect 46924 18332 46964 18451
rect 47020 18450 47060 18535
rect 47404 18450 47444 18535
rect 47500 18425 47540 18544
rect 47596 18584 47636 18712
rect 47499 18416 47541 18425
rect 47499 18376 47500 18416
rect 47540 18376 47541 18416
rect 47499 18367 47541 18376
rect 47020 18332 47060 18341
rect 46924 18292 47020 18332
rect 47020 18283 47060 18292
rect 46827 17324 46869 17333
rect 46827 17284 46828 17324
rect 46868 17284 46869 17324
rect 46827 17275 46869 17284
rect 47596 17240 47636 18544
rect 47691 18584 47733 18593
rect 47691 18544 47692 18584
rect 47732 18544 47733 18584
rect 47691 18535 47733 18544
rect 47692 18450 47732 18535
rect 45812 17116 46100 17156
rect 46540 17200 46676 17240
rect 47404 17200 47636 17240
rect 45676 17072 45716 17083
rect 45676 16997 45716 17032
rect 45675 16988 45717 16997
rect 45675 16948 45676 16988
rect 45716 16948 45717 16988
rect 45675 16939 45717 16948
rect 45676 16484 45716 16493
rect 45772 16484 45812 17116
rect 46252 17072 46292 17081
rect 45867 16820 45909 16829
rect 45867 16780 45868 16820
rect 45908 16780 45909 16820
rect 45867 16771 45909 16780
rect 46060 16820 46100 16829
rect 46100 16780 46196 16820
rect 46060 16771 46100 16780
rect 45716 16444 45812 16484
rect 45676 16435 45716 16444
rect 45868 16232 45908 16771
rect 45963 16568 46005 16577
rect 45963 16528 45964 16568
rect 46004 16528 46005 16568
rect 45963 16519 46005 16528
rect 45964 16484 46004 16519
rect 45964 16433 46004 16444
rect 46156 16400 46196 16780
rect 46252 16577 46292 17032
rect 46251 16568 46293 16577
rect 46251 16528 46252 16568
rect 46292 16528 46293 16568
rect 46251 16519 46293 16528
rect 46156 16360 46388 16400
rect 45964 16232 46004 16241
rect 46156 16232 46196 16241
rect 45868 16192 45964 16232
rect 45964 16183 46004 16192
rect 46060 16192 46156 16232
rect 45579 16148 45621 16157
rect 45579 16108 45580 16148
rect 45620 16108 45621 16148
rect 45579 16099 45621 16108
rect 45483 16064 45525 16073
rect 45483 16024 45484 16064
rect 45524 16024 45525 16064
rect 45483 16015 45525 16024
rect 45676 16064 45716 16073
rect 45483 15728 45525 15737
rect 45483 15688 45484 15728
rect 45524 15688 45525 15728
rect 45483 15679 45525 15688
rect 45388 15560 45428 15569
rect 45388 15308 45428 15520
rect 45484 15560 45524 15679
rect 45579 15644 45621 15653
rect 45579 15604 45580 15644
rect 45620 15604 45621 15644
rect 45579 15595 45621 15604
rect 45484 15511 45524 15520
rect 45580 15560 45620 15595
rect 45580 15509 45620 15520
rect 45676 15560 45716 16024
rect 45963 15896 46005 15905
rect 45963 15856 45964 15896
rect 46004 15856 46005 15896
rect 45963 15847 46005 15856
rect 45964 15728 46004 15847
rect 45964 15679 46004 15688
rect 46060 15569 46100 16192
rect 46156 16183 46196 16192
rect 46251 16232 46293 16241
rect 46251 16192 46252 16232
rect 46292 16192 46293 16232
rect 46251 16183 46293 16192
rect 46252 16098 46292 16183
rect 46251 15644 46293 15653
rect 46251 15604 46252 15644
rect 46292 15604 46293 15644
rect 46251 15595 46293 15604
rect 45676 15511 45716 15520
rect 45868 15560 45908 15569
rect 45868 15308 45908 15520
rect 46059 15560 46101 15569
rect 46059 15520 46060 15560
rect 46100 15520 46101 15560
rect 46059 15511 46101 15520
rect 46156 15560 46196 15569
rect 46060 15426 46100 15511
rect 45388 15268 45908 15308
rect 46156 14981 46196 15520
rect 46252 15308 46292 15595
rect 46348 15560 46388 16360
rect 46540 16316 46580 17200
rect 46636 17072 46676 17081
rect 46676 17032 46868 17072
rect 46636 17023 46676 17032
rect 46828 16400 46868 17032
rect 47211 16904 47253 16913
rect 47211 16864 47212 16904
rect 47252 16864 47253 16904
rect 47211 16855 47253 16864
rect 46828 16351 46868 16360
rect 46636 16316 46676 16325
rect 46540 16276 46636 16316
rect 46636 16267 46676 16276
rect 46444 16064 46484 16073
rect 46484 16024 46580 16064
rect 46444 16015 46484 16024
rect 46348 15511 46388 15520
rect 46443 15560 46485 15569
rect 46443 15520 46444 15560
rect 46484 15520 46485 15560
rect 46443 15511 46485 15520
rect 46540 15560 46580 16024
rect 47212 15728 47252 16855
rect 47164 15688 47252 15728
rect 47164 15644 47204 15688
rect 47404 15653 47444 17200
rect 47500 17072 47540 17081
rect 47788 17072 47828 19216
rect 48075 18668 48117 18677
rect 48075 18628 48076 18668
rect 48116 18628 48117 18668
rect 48075 18619 48117 18628
rect 47980 18584 48020 18593
rect 47980 18509 48020 18544
rect 48076 18534 48116 18619
rect 48172 18584 48212 18593
rect 47979 18500 48021 18509
rect 47979 18460 47980 18500
rect 48020 18460 48021 18500
rect 47979 18451 48021 18460
rect 47980 17417 48020 18451
rect 48172 18416 48212 18544
rect 48364 18416 48404 18425
rect 48172 18376 48364 18416
rect 48364 18367 48404 18376
rect 48460 18341 48500 19636
rect 49132 19508 49172 19804
rect 48844 19468 49172 19508
rect 48748 19088 48788 19097
rect 48652 19048 48748 19088
rect 48652 18668 48692 19048
rect 48748 19039 48788 19048
rect 48652 18593 48692 18628
rect 48651 18584 48693 18593
rect 48651 18544 48652 18584
rect 48692 18544 48693 18584
rect 48651 18535 48693 18544
rect 48748 18584 48788 18593
rect 48459 18332 48501 18341
rect 48459 18292 48460 18332
rect 48500 18292 48501 18332
rect 48459 18283 48501 18292
rect 48267 18164 48309 18173
rect 48267 18124 48268 18164
rect 48308 18124 48309 18164
rect 48267 18115 48309 18124
rect 48268 17828 48308 18115
rect 48459 17912 48501 17921
rect 48459 17872 48460 17912
rect 48500 17872 48501 17912
rect 48459 17863 48501 17872
rect 48268 17779 48308 17788
rect 48460 17778 48500 17863
rect 48652 17744 48692 18535
rect 48748 18425 48788 18544
rect 48844 18509 48884 19468
rect 49036 19256 49076 19265
rect 48939 18920 48981 18929
rect 48939 18880 48940 18920
rect 48980 18880 48981 18920
rect 48939 18871 48981 18880
rect 48940 18593 48980 18871
rect 49036 18761 49076 19216
rect 49228 19256 49268 19265
rect 49131 19172 49173 19181
rect 49131 19132 49132 19172
rect 49172 19132 49173 19172
rect 49131 19123 49173 19132
rect 49132 19038 49172 19123
rect 49228 18761 49268 19216
rect 49324 19256 49364 19265
rect 49035 18752 49077 18761
rect 49035 18712 49036 18752
rect 49076 18712 49077 18752
rect 49035 18703 49077 18712
rect 49227 18752 49269 18761
rect 49227 18712 49228 18752
rect 49268 18712 49269 18752
rect 49324 18752 49364 19216
rect 49996 19256 50036 19888
rect 50092 19879 50132 19888
rect 49996 19207 50036 19216
rect 50860 19256 50900 20719
rect 51532 20634 51572 20719
rect 51627 20012 51669 20021
rect 51627 19972 51628 20012
rect 51668 19972 51669 20012
rect 51627 19963 51669 19972
rect 50860 19207 50900 19216
rect 49611 19172 49653 19181
rect 49611 19132 49612 19172
rect 49652 19132 49653 19172
rect 49611 19123 49653 19132
rect 49612 19038 49652 19123
rect 50859 18836 50901 18845
rect 50859 18796 50860 18836
rect 50900 18796 50901 18836
rect 50859 18787 50901 18796
rect 49324 18712 49460 18752
rect 49227 18703 49269 18712
rect 49420 18668 49460 18712
rect 49420 18619 49460 18628
rect 48939 18584 48981 18593
rect 48939 18544 48940 18584
rect 48980 18544 48981 18584
rect 48939 18535 48981 18544
rect 49036 18584 49076 18593
rect 49324 18584 49364 18593
rect 49076 18544 49268 18584
rect 49036 18535 49076 18544
rect 48843 18500 48885 18509
rect 48843 18460 48844 18500
rect 48884 18460 48885 18500
rect 48843 18451 48885 18460
rect 48747 18416 48789 18425
rect 48747 18376 48748 18416
rect 48788 18376 48789 18416
rect 48747 18367 48789 18376
rect 48939 17912 48981 17921
rect 48939 17872 48940 17912
rect 48980 17872 48981 17912
rect 48939 17863 48981 17872
rect 48652 17695 48692 17704
rect 48748 17744 48788 17753
rect 48748 17585 48788 17704
rect 48940 17744 48980 17863
rect 48980 17704 49076 17744
rect 48940 17695 48980 17704
rect 48747 17576 48789 17585
rect 48747 17536 48748 17576
rect 48788 17536 48789 17576
rect 48747 17527 48789 17536
rect 48844 17576 48884 17585
rect 47979 17408 48021 17417
rect 47979 17368 47980 17408
rect 48020 17368 48021 17408
rect 47979 17359 48021 17368
rect 48844 17333 48884 17536
rect 48939 17408 48981 17417
rect 48939 17368 48940 17408
rect 48980 17368 48981 17408
rect 48939 17359 48981 17368
rect 48843 17324 48885 17333
rect 48843 17284 48844 17324
rect 48884 17284 48885 17324
rect 48843 17275 48885 17284
rect 48267 17240 48309 17249
rect 48267 17200 48268 17240
rect 48308 17200 48309 17240
rect 48267 17191 48309 17200
rect 47540 17032 47828 17072
rect 47500 17023 47540 17032
rect 48268 16913 48308 17191
rect 48651 16988 48693 16997
rect 48651 16948 48652 16988
rect 48692 16948 48693 16988
rect 48651 16939 48693 16948
rect 48267 16904 48309 16913
rect 48267 16864 48268 16904
rect 48308 16864 48309 16904
rect 48267 16855 48309 16864
rect 48652 16854 48692 16939
rect 48651 16232 48693 16241
rect 48651 16192 48652 16232
rect 48692 16192 48693 16232
rect 48651 16183 48693 16192
rect 48652 16098 48692 16183
rect 47116 15604 47204 15644
rect 47403 15644 47445 15653
rect 47403 15604 47404 15644
rect 47444 15604 47445 15644
rect 46444 15426 46484 15511
rect 46252 15268 46484 15308
rect 45579 14972 45621 14981
rect 45579 14932 45580 14972
rect 45620 14932 45621 14972
rect 45579 14923 45621 14932
rect 46155 14972 46197 14981
rect 46155 14932 46156 14972
rect 46196 14932 46197 14972
rect 46155 14923 46197 14932
rect 45580 14838 45620 14923
rect 45771 14804 45813 14813
rect 45292 14764 45524 14804
rect 45484 14720 45524 14764
rect 45771 14764 45772 14804
rect 45812 14764 45813 14804
rect 45771 14755 45813 14764
rect 45580 14720 45620 14729
rect 45484 14680 45580 14720
rect 45044 14008 45140 14048
rect 45004 13999 45044 14008
rect 45483 13460 45525 13469
rect 45483 13420 45484 13460
rect 45524 13420 45525 13460
rect 45483 13411 45525 13420
rect 45484 13326 45524 13411
rect 44811 12704 44853 12713
rect 44811 12664 44812 12704
rect 44852 12664 44853 12704
rect 44811 12655 44853 12664
rect 45484 12536 45524 12545
rect 44715 12200 44757 12209
rect 44715 12160 44716 12200
rect 44756 12160 44757 12200
rect 44715 12151 44757 12160
rect 44619 12032 44661 12041
rect 44619 11992 44620 12032
rect 44660 11992 44661 12032
rect 44619 11983 44661 11992
rect 44716 11948 44756 12151
rect 45484 11957 45524 12496
rect 45580 12293 45620 14680
rect 45772 14720 45812 14755
rect 45772 14669 45812 14680
rect 45867 14720 45909 14729
rect 45867 14680 45868 14720
rect 45908 14680 45909 14720
rect 45867 14671 45909 14680
rect 46252 14720 46292 14729
rect 45868 14586 45908 14671
rect 46252 14645 46292 14680
rect 46347 14720 46389 14729
rect 46347 14680 46348 14720
rect 46388 14680 46389 14720
rect 46347 14671 46389 14680
rect 46251 14636 46293 14645
rect 46251 14596 46252 14636
rect 46292 14596 46293 14636
rect 46251 14587 46293 14596
rect 46059 14384 46101 14393
rect 46059 14344 46060 14384
rect 46100 14344 46101 14384
rect 46059 14335 46101 14344
rect 45867 14132 45909 14141
rect 45867 14092 45868 14132
rect 45908 14092 45909 14132
rect 45867 14083 45909 14092
rect 45868 14048 45908 14083
rect 45868 13997 45908 14008
rect 46060 13385 46100 14335
rect 46252 14141 46292 14587
rect 46251 14132 46293 14141
rect 46251 14092 46252 14132
rect 46292 14092 46293 14132
rect 46251 14083 46293 14092
rect 46155 14048 46197 14057
rect 46155 14008 46156 14048
rect 46196 14008 46197 14048
rect 46155 13999 46197 14008
rect 46059 13376 46101 13385
rect 46059 13336 46060 13376
rect 46100 13336 46101 13376
rect 46059 13327 46101 13336
rect 46156 13208 46196 13999
rect 46156 13159 46196 13168
rect 46252 13049 46292 14083
rect 46348 13124 46388 14671
rect 46348 13084 46391 13124
rect 46251 13040 46293 13049
rect 46351 13040 46391 13084
rect 46251 13000 46252 13040
rect 46292 13000 46293 13040
rect 46251 12991 46293 13000
rect 46348 13000 46391 13040
rect 45868 12536 45908 12545
rect 45579 12284 45621 12293
rect 45579 12244 45580 12284
rect 45620 12244 45621 12284
rect 45579 12235 45621 12244
rect 44716 11899 44756 11908
rect 45483 11948 45525 11957
rect 45483 11908 45484 11948
rect 45524 11908 45525 11948
rect 45483 11899 45525 11908
rect 44523 11864 44565 11873
rect 44523 11824 44524 11864
rect 44564 11824 44565 11864
rect 44523 11815 44565 11824
rect 44907 11864 44949 11873
rect 44907 11824 44908 11864
rect 44948 11824 44949 11864
rect 45868 11864 45908 12496
rect 45964 11864 46004 11873
rect 45868 11824 45964 11864
rect 44907 11815 44949 11824
rect 45964 11815 46004 11824
rect 44524 11024 44564 11815
rect 44908 11730 44948 11815
rect 45387 11696 45429 11705
rect 45387 11656 45388 11696
rect 45428 11656 45429 11696
rect 45387 11647 45429 11656
rect 46348 11696 46388 13000
rect 46348 11647 46388 11656
rect 46444 11696 46484 15268
rect 46540 14393 46580 15520
rect 46924 15560 46964 15569
rect 47116 15560 47156 15604
rect 47403 15595 47445 15604
rect 48075 15644 48117 15653
rect 48075 15604 48076 15644
rect 48116 15604 48117 15644
rect 48075 15595 48117 15604
rect 46964 15520 47156 15560
rect 47308 15560 47348 15569
rect 46924 14561 46964 15520
rect 47212 15518 47252 15527
rect 47212 15401 47252 15478
rect 47211 15392 47253 15401
rect 47211 15352 47212 15392
rect 47252 15352 47253 15392
rect 47211 15343 47253 15352
rect 47308 14729 47348 15520
rect 47788 15560 47828 15569
rect 47788 15401 47828 15520
rect 47979 15560 48021 15569
rect 47979 15520 47980 15560
rect 48020 15520 48021 15560
rect 47979 15511 48021 15520
rect 47980 15426 48020 15511
rect 47787 15392 47829 15401
rect 47787 15352 47788 15392
rect 47828 15352 47829 15392
rect 47787 15343 47829 15352
rect 47596 15308 47636 15317
rect 47307 14720 47349 14729
rect 47307 14680 47308 14720
rect 47348 14680 47349 14720
rect 47307 14671 47349 14680
rect 47404 14720 47444 14729
rect 46923 14552 46965 14561
rect 46923 14512 46924 14552
rect 46964 14512 46965 14552
rect 46923 14503 46965 14512
rect 46539 14384 46581 14393
rect 46539 14344 46540 14384
rect 46580 14344 46581 14384
rect 46539 14335 46581 14344
rect 46539 14048 46581 14057
rect 47308 14048 47348 14671
rect 47404 14393 47444 14680
rect 47596 14720 47636 15268
rect 47596 14671 47636 14680
rect 47884 15308 47924 15317
rect 47500 14636 47540 14645
rect 47403 14384 47445 14393
rect 47403 14344 47404 14384
rect 47444 14344 47445 14384
rect 47403 14335 47445 14344
rect 47500 14057 47540 14596
rect 47595 14132 47637 14141
rect 47595 14092 47596 14132
rect 47636 14092 47637 14132
rect 47595 14083 47637 14092
rect 47692 14132 47732 14141
rect 46539 14008 46540 14048
rect 46580 14008 46581 14048
rect 46539 13999 46581 14008
rect 47020 14008 47348 14048
rect 47499 14048 47541 14057
rect 47499 14008 47500 14048
rect 47540 14008 47541 14048
rect 46540 13544 46580 13999
rect 47020 13964 47060 14008
rect 47499 13999 47541 14008
rect 47596 14048 47636 14083
rect 47596 13997 47636 14008
rect 47020 13915 47060 13924
rect 47692 13880 47732 14092
rect 47788 14057 47828 14142
rect 47787 14048 47829 14057
rect 47787 14008 47788 14048
rect 47828 14008 47829 14048
rect 47787 13999 47829 14008
rect 47884 14048 47924 15268
rect 47884 13999 47924 14008
rect 47980 14636 48020 14645
rect 47980 13880 48020 14596
rect 47692 13840 48020 13880
rect 48076 13796 48116 15595
rect 48460 15392 48500 15401
rect 48364 15352 48460 15392
rect 48364 14720 48404 15352
rect 48460 15343 48500 15352
rect 48940 15317 48980 17359
rect 49036 16904 49076 17704
rect 49131 17324 49173 17333
rect 49131 17284 49132 17324
rect 49172 17284 49173 17324
rect 49131 17275 49173 17284
rect 49132 17072 49172 17275
rect 49228 17249 49268 18544
rect 49324 18257 49364 18544
rect 49516 18584 49556 18595
rect 49900 18593 49940 18624
rect 49516 18509 49556 18544
rect 49899 18584 49941 18593
rect 49899 18544 49900 18584
rect 49940 18544 49941 18584
rect 49899 18535 49941 18544
rect 49515 18500 49557 18509
rect 49515 18460 49516 18500
rect 49556 18460 49557 18500
rect 49515 18451 49557 18460
rect 49900 18500 49940 18535
rect 49900 18341 49940 18460
rect 50572 18500 50612 18509
rect 49419 18332 49461 18341
rect 49419 18292 49420 18332
rect 49460 18292 49461 18332
rect 49419 18283 49461 18292
rect 49899 18332 49941 18341
rect 50092 18332 50132 18341
rect 49899 18292 49900 18332
rect 49940 18292 49941 18332
rect 49899 18283 49941 18292
rect 49996 18292 50092 18332
rect 49323 18248 49365 18257
rect 49323 18208 49324 18248
rect 49364 18208 49365 18248
rect 49323 18199 49365 18208
rect 49420 17921 49460 18283
rect 49419 17912 49461 17921
rect 49419 17872 49420 17912
rect 49460 17872 49461 17912
rect 49419 17863 49461 17872
rect 49516 17872 49940 17912
rect 49420 17828 49460 17863
rect 49420 17777 49460 17788
rect 49516 17660 49556 17872
rect 49900 17758 49940 17872
rect 49324 17620 49556 17660
rect 49804 17744 49844 17753
rect 49900 17709 49940 17718
rect 49804 17660 49844 17704
rect 49804 17620 49940 17660
rect 49227 17240 49269 17249
rect 49227 17200 49228 17240
rect 49268 17200 49269 17240
rect 49227 17191 49269 17200
rect 49132 17023 49172 17032
rect 49228 17072 49268 17081
rect 49324 17072 49364 17620
rect 49612 17576 49652 17585
rect 49652 17536 49844 17576
rect 49612 17527 49652 17536
rect 49268 17032 49364 17072
rect 49420 17072 49460 17081
rect 49460 17032 49748 17072
rect 49228 16913 49268 17032
rect 49420 17023 49460 17032
rect 49227 16904 49269 16913
rect 49036 16864 49172 16904
rect 49036 16232 49076 16241
rect 49036 15392 49076 16192
rect 49132 15653 49172 16864
rect 49227 16864 49228 16904
rect 49268 16864 49269 16904
rect 49227 16855 49269 16864
rect 49323 16820 49365 16829
rect 49323 16780 49324 16820
rect 49364 16780 49365 16820
rect 49323 16771 49365 16780
rect 49420 16820 49460 16829
rect 49131 15644 49173 15653
rect 49131 15604 49132 15644
rect 49172 15604 49173 15644
rect 49131 15595 49173 15604
rect 49132 15392 49172 15401
rect 49036 15352 49132 15392
rect 49132 15343 49172 15352
rect 48939 15308 48981 15317
rect 48939 15268 48940 15308
rect 48980 15268 48981 15308
rect 48939 15259 48981 15268
rect 48364 14671 48404 14680
rect 49228 14720 49268 14731
rect 49228 14645 49268 14680
rect 49227 14636 49269 14645
rect 49227 14596 49228 14636
rect 49268 14596 49269 14636
rect 49227 14587 49269 14596
rect 48363 14552 48405 14561
rect 48363 14512 48364 14552
rect 48404 14512 48405 14552
rect 48363 14503 48405 14512
rect 47980 13756 48116 13796
rect 46540 13504 46868 13544
rect 46635 13040 46677 13049
rect 46635 13000 46636 13040
rect 46676 13000 46772 13040
rect 46635 12991 46677 13000
rect 46636 12906 46676 12991
rect 46732 12536 46772 13000
rect 46732 12487 46772 12496
rect 46828 12461 46868 13504
rect 47020 13504 47348 13544
rect 47020 13208 47060 13504
rect 47308 13460 47348 13504
rect 47308 13411 47348 13420
rect 47500 13301 47540 13317
rect 47499 13292 47541 13301
rect 47499 13252 47500 13292
rect 47540 13252 47541 13292
rect 47499 13243 47541 13252
rect 47500 13222 47540 13243
rect 46924 13168 47060 13208
rect 47308 13208 47348 13217
rect 47500 13173 47540 13182
rect 47596 13208 47636 13217
rect 47884 13208 47924 13217
rect 46827 12452 46869 12461
rect 46827 12412 46828 12452
rect 46868 12412 46869 12452
rect 46827 12403 46869 12412
rect 46827 12032 46869 12041
rect 46827 11992 46828 12032
rect 46868 11992 46869 12032
rect 46827 11983 46869 11992
rect 46828 11948 46868 11983
rect 46828 11897 46868 11908
rect 46539 11780 46581 11789
rect 46539 11740 46540 11780
rect 46580 11740 46581 11780
rect 46539 11731 46581 11740
rect 46444 11647 46484 11656
rect 46540 11696 46580 11731
rect 46924 11705 46964 13168
rect 47308 13124 47348 13168
rect 47636 13168 47884 13208
rect 47596 13159 47636 13168
rect 47308 13084 47492 13124
rect 47452 13040 47492 13084
rect 47452 13000 47540 13040
rect 47500 12881 47540 13000
rect 47499 12872 47541 12881
rect 47499 12832 47500 12872
rect 47540 12832 47541 12872
rect 47499 12823 47541 12832
rect 47884 12713 47924 13168
rect 47980 13208 48020 13756
rect 48075 13460 48117 13469
rect 48075 13420 48076 13460
rect 48116 13420 48117 13460
rect 48075 13411 48117 13420
rect 48076 13250 48116 13411
rect 48076 13201 48116 13210
rect 47980 13159 48020 13168
rect 48172 13040 48212 13049
rect 48172 12980 48212 13000
rect 48076 12940 48212 12980
rect 47883 12704 47925 12713
rect 47883 12664 47884 12704
rect 47924 12664 47925 12704
rect 47883 12655 47925 12664
rect 47884 12570 47924 12655
rect 47019 12452 47061 12461
rect 47019 12412 47020 12452
rect 47060 12412 47061 12452
rect 47019 12403 47061 12412
rect 44524 10975 44564 10984
rect 45388 11024 45428 11647
rect 46540 11645 46580 11656
rect 46636 11696 46676 11705
rect 46828 11696 46868 11705
rect 46676 11656 46828 11696
rect 46636 11647 46676 11656
rect 46828 11647 46868 11656
rect 46923 11696 46965 11705
rect 46923 11656 46924 11696
rect 46964 11656 46965 11696
rect 46923 11647 46965 11656
rect 47020 11696 47060 12403
rect 47020 11647 47060 11656
rect 47115 11696 47157 11705
rect 47115 11656 47116 11696
rect 47156 11656 47157 11696
rect 48076 11696 48116 12940
rect 48172 12536 48212 12545
rect 48364 12536 48404 14503
rect 48651 14384 48693 14393
rect 48651 14344 48652 14384
rect 48692 14344 48693 14384
rect 48651 14335 48693 14344
rect 48459 13376 48501 13385
rect 48459 13336 48460 13376
rect 48500 13336 48501 13376
rect 48459 13327 48501 13336
rect 48460 13049 48500 13327
rect 48652 13208 48692 14335
rect 49324 14141 49364 16771
rect 49420 16241 49460 16780
rect 49419 16232 49461 16241
rect 49419 16192 49420 16232
rect 49460 16192 49461 16232
rect 49419 16183 49461 16192
rect 49708 15728 49748 17032
rect 49708 15679 49748 15688
rect 49804 15560 49844 17536
rect 49900 17165 49940 17620
rect 49899 17156 49941 17165
rect 49899 17116 49900 17156
rect 49940 17116 49941 17156
rect 49899 17107 49941 17116
rect 49900 16988 49940 16997
rect 49900 16829 49940 16948
rect 49899 16820 49941 16829
rect 49899 16780 49900 16820
rect 49940 16780 49941 16820
rect 49899 16771 49941 16780
rect 49900 16232 49940 16241
rect 49900 15905 49940 16192
rect 49899 15896 49941 15905
rect 49899 15856 49900 15896
rect 49940 15856 49941 15896
rect 49899 15847 49941 15856
rect 49996 15728 50036 18292
rect 50092 18283 50132 18292
rect 50380 18332 50420 18341
rect 50092 17912 50132 17921
rect 50132 17872 50324 17912
rect 50092 17863 50132 17872
rect 50091 17744 50133 17753
rect 50091 17704 50092 17744
rect 50132 17704 50133 17744
rect 50091 17695 50133 17704
rect 50284 17744 50324 17872
rect 50380 17753 50420 18292
rect 50572 18173 50612 18460
rect 50764 18416 50804 18425
rect 50571 18164 50613 18173
rect 50571 18124 50572 18164
rect 50612 18124 50613 18164
rect 50571 18115 50613 18124
rect 50571 17912 50613 17921
rect 50571 17872 50572 17912
rect 50612 17872 50613 17912
rect 50571 17863 50613 17872
rect 50475 17828 50517 17837
rect 50475 17788 50476 17828
rect 50516 17788 50517 17828
rect 50475 17779 50517 17788
rect 50284 17695 50324 17704
rect 50379 17744 50421 17753
rect 50379 17704 50380 17744
rect 50420 17704 50421 17744
rect 50379 17695 50421 17704
rect 50092 17610 50132 17695
rect 50380 17072 50420 17081
rect 50092 16820 50132 16829
rect 50380 16820 50420 17032
rect 50132 16780 50420 16820
rect 50092 16771 50132 16780
rect 49925 15688 50228 15728
rect 49925 15644 49965 15688
rect 49708 15520 49804 15560
rect 49035 14132 49077 14141
rect 49035 14092 49036 14132
rect 49076 14092 49077 14132
rect 49035 14083 49077 14092
rect 49323 14132 49365 14141
rect 49323 14092 49324 14132
rect 49364 14092 49365 14132
rect 49323 14083 49365 14092
rect 48652 13159 48692 13168
rect 48844 13208 48884 13217
rect 48748 13124 48788 13133
rect 48459 13040 48501 13049
rect 48459 13000 48460 13040
rect 48500 13000 48501 13040
rect 48459 12991 48501 13000
rect 48459 12788 48501 12797
rect 48459 12748 48460 12788
rect 48500 12748 48501 12788
rect 48459 12739 48501 12748
rect 48212 12496 48404 12536
rect 48460 12536 48500 12739
rect 48748 12713 48788 13084
rect 48555 12704 48597 12713
rect 48555 12664 48556 12704
rect 48596 12664 48597 12704
rect 48555 12655 48597 12664
rect 48747 12704 48789 12713
rect 48747 12664 48748 12704
rect 48788 12664 48789 12704
rect 48747 12655 48789 12664
rect 48556 12620 48596 12655
rect 48556 12569 48596 12580
rect 48172 12487 48212 12496
rect 48460 12487 48500 12496
rect 48844 12368 48884 13168
rect 49036 12536 49076 14083
rect 49515 13292 49557 13301
rect 49515 13252 49516 13292
rect 49556 13252 49557 13292
rect 49515 13243 49557 13252
rect 49131 13124 49173 13133
rect 49131 13084 49132 13124
rect 49172 13084 49173 13124
rect 49131 13075 49173 13084
rect 49419 13124 49461 13133
rect 49419 13084 49420 13124
rect 49460 13084 49461 13124
rect 49419 13075 49461 13084
rect 49132 12704 49172 13075
rect 49420 12990 49460 13075
rect 49132 12655 49172 12664
rect 49227 12704 49269 12713
rect 49227 12664 49228 12704
rect 49268 12664 49269 12704
rect 49227 12655 49269 12664
rect 49036 12487 49076 12496
rect 49228 12536 49268 12655
rect 48844 12319 48884 12328
rect 48267 11948 48309 11957
rect 48267 11908 48268 11948
rect 48308 11908 48309 11948
rect 48267 11899 48309 11908
rect 48268 11814 48308 11899
rect 49132 11873 49172 11958
rect 48555 11864 48597 11873
rect 48555 11824 48556 11864
rect 48596 11824 48597 11864
rect 48555 11815 48597 11824
rect 49131 11864 49173 11873
rect 49131 11824 49132 11864
rect 49172 11824 49173 11864
rect 49131 11815 49173 11824
rect 48268 11696 48308 11705
rect 48076 11656 48268 11696
rect 47115 11647 47157 11656
rect 48268 11647 48308 11656
rect 48459 11696 48501 11705
rect 48459 11656 48460 11696
rect 48500 11656 48501 11696
rect 48459 11647 48501 11656
rect 48556 11696 48596 11815
rect 49228 11705 49268 12496
rect 49323 12536 49365 12545
rect 49323 12496 49324 12536
rect 49364 12496 49365 12536
rect 49323 12487 49365 12496
rect 49516 12536 49556 13243
rect 49708 12881 49748 15520
rect 49804 15511 49844 15520
rect 49900 15604 49965 15644
rect 49900 15560 49940 15604
rect 49900 15511 49940 15520
rect 49995 15560 50037 15569
rect 49995 15520 49996 15560
rect 50036 15520 50037 15560
rect 49995 15511 50037 15520
rect 49996 15426 50036 15511
rect 49995 15308 50037 15317
rect 49995 15268 49996 15308
rect 50036 15268 50037 15308
rect 49995 15259 50037 15268
rect 49804 13208 49844 13217
rect 49804 12980 49844 13168
rect 49804 12940 49940 12980
rect 49707 12872 49749 12881
rect 49707 12832 49708 12872
rect 49748 12832 49749 12872
rect 49707 12823 49749 12832
rect 49707 12704 49749 12713
rect 49707 12664 49708 12704
rect 49748 12664 49749 12704
rect 49707 12655 49749 12664
rect 49324 12402 49364 12487
rect 49516 12284 49556 12496
rect 49611 12536 49653 12545
rect 49611 12496 49612 12536
rect 49652 12496 49653 12536
rect 49611 12487 49653 12496
rect 49708 12536 49748 12655
rect 49708 12487 49748 12496
rect 49612 12402 49652 12487
rect 49900 12368 49940 12940
rect 49900 12319 49940 12328
rect 49324 12244 49556 12284
rect 49611 12284 49653 12293
rect 49611 12244 49612 12284
rect 49652 12244 49653 12284
rect 48556 11647 48596 11656
rect 49132 11696 49172 11705
rect 47116 11562 47156 11647
rect 48460 11562 48500 11647
rect 49132 11537 49172 11656
rect 49227 11696 49269 11705
rect 49227 11656 49228 11696
rect 49268 11656 49269 11696
rect 49227 11647 49269 11656
rect 49324 11696 49364 12244
rect 49611 12235 49653 12244
rect 49612 11780 49652 12235
rect 49612 11731 49652 11740
rect 49804 11864 49844 11873
rect 49324 11647 49364 11656
rect 49419 11696 49461 11705
rect 49419 11656 49420 11696
rect 49460 11656 49461 11696
rect 49419 11647 49461 11656
rect 49420 11562 49460 11647
rect 49804 11537 49844 11824
rect 49131 11528 49173 11537
rect 49131 11488 49132 11528
rect 49172 11488 49173 11528
rect 49131 11479 49173 11488
rect 49803 11528 49845 11537
rect 49803 11488 49804 11528
rect 49844 11488 49845 11528
rect 49803 11479 49845 11488
rect 46251 11276 46293 11285
rect 46251 11236 46252 11276
rect 46292 11236 46293 11276
rect 46251 11227 46293 11236
rect 45388 10975 45428 10984
rect 46252 10277 46292 11227
rect 46539 11192 46581 11201
rect 46539 11152 46540 11192
rect 46580 11152 46581 11192
rect 46539 11143 46581 11152
rect 46732 11152 47060 11192
rect 46540 10865 46580 11143
rect 46539 10856 46581 10865
rect 46539 10816 46540 10856
rect 46580 10816 46581 10856
rect 46539 10807 46581 10816
rect 46540 10722 46580 10807
rect 46732 10436 46772 11152
rect 47020 11108 47060 11152
rect 47020 11059 47060 11068
rect 48075 11108 48117 11117
rect 48075 11068 48076 11108
rect 48116 11068 48117 11108
rect 48075 11059 48117 11068
rect 46924 11024 46964 11033
rect 46540 10396 46772 10436
rect 46827 10436 46869 10445
rect 46827 10396 46828 10436
rect 46868 10396 46869 10436
rect 46251 10268 46293 10277
rect 44428 10228 44564 10268
rect 44332 10135 44372 10144
rect 44524 10184 44564 10228
rect 46251 10228 46252 10268
rect 46292 10228 46293 10268
rect 46251 10219 46293 10228
rect 43659 10100 43701 10109
rect 43659 10060 43660 10100
rect 43700 10060 43701 10100
rect 43659 10051 43701 10060
rect 43852 10100 43892 10109
rect 43275 9932 43317 9941
rect 43275 9892 43276 9932
rect 43316 9892 43317 9932
rect 43275 9883 43317 9892
rect 43083 9680 43125 9689
rect 43083 9640 43084 9680
rect 43124 9640 43125 9680
rect 43083 9631 43125 9640
rect 42987 9596 43029 9605
rect 42987 9556 42988 9596
rect 43028 9556 43029 9596
rect 42987 9547 43029 9556
rect 42796 9463 42836 9472
rect 42891 9512 42933 9521
rect 42891 9472 42892 9512
rect 42932 9472 42933 9512
rect 42891 9463 42933 9472
rect 42700 9378 42740 9463
rect 42892 9378 42932 9463
rect 41972 9304 42164 9344
rect 41932 9295 41972 9304
rect 42411 9260 42453 9269
rect 42411 9220 42412 9260
rect 42452 9220 42453 9260
rect 42411 9211 42453 9220
rect 42412 9126 42452 9211
rect 41835 8756 41877 8765
rect 41835 8716 41836 8756
rect 41876 8716 41877 8756
rect 41835 8707 41877 8716
rect 42795 8756 42837 8765
rect 42795 8716 42796 8756
rect 42836 8716 42837 8756
rect 42795 8707 42837 8716
rect 41931 8672 41973 8681
rect 41931 8632 41932 8672
rect 41972 8632 41973 8672
rect 41931 8623 41973 8632
rect 42796 8672 42836 8707
rect 41548 8539 41588 8548
rect 41932 8538 41972 8623
rect 42796 8621 42836 8632
rect 7659 8504 7701 8513
rect 7659 8464 7660 8504
rect 7700 8464 7701 8504
rect 7659 8455 7701 8464
rect 7468 8119 7508 8128
rect 6316 8000 6356 8009
rect 6028 7960 6316 8000
rect 6316 7951 6356 7960
rect 6411 8000 6453 8009
rect 6411 7960 6412 8000
rect 6452 7960 6453 8000
rect 6411 7951 6453 7960
rect 6316 6488 6356 6497
rect 6220 6448 6316 6488
rect 6220 5657 6260 6448
rect 6316 6439 6356 6448
rect 6316 5909 6356 5994
rect 6315 5900 6357 5909
rect 6315 5860 6316 5900
rect 6356 5860 6357 5900
rect 6315 5851 6357 5860
rect 6028 5648 6068 5657
rect 5932 5608 6028 5648
rect 5932 5153 5972 5608
rect 6028 5599 6068 5608
rect 6124 5648 6164 5657
rect 6124 5237 6164 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6316 5648 6356 5657
rect 6412 5648 6452 7951
rect 7467 7748 7509 7757
rect 7467 7708 7468 7748
rect 7508 7708 7509 7748
rect 7467 7699 7509 7708
rect 7468 7614 7508 7699
rect 7468 6656 7508 6667
rect 7468 6581 7508 6616
rect 7467 6572 7509 6581
rect 7467 6532 7468 6572
rect 7508 6532 7509 6572
rect 7467 6523 7509 6532
rect 7468 6245 7508 6523
rect 7467 6236 7509 6245
rect 7467 6196 7468 6236
rect 7508 6196 7509 6236
rect 7467 6187 7509 6196
rect 6356 5608 6452 5648
rect 6123 5228 6165 5237
rect 6123 5188 6124 5228
rect 6164 5188 6165 5228
rect 6123 5179 6165 5188
rect 5931 5144 5973 5153
rect 5931 5104 5932 5144
rect 5972 5104 5973 5144
rect 5931 5095 5973 5104
rect 5836 4936 6068 4976
rect 5548 4808 5588 4817
rect 5932 4808 5972 4817
rect 5452 4768 5548 4808
rect 5548 4759 5588 4768
rect 5740 4768 5932 4808
rect 5068 4304 5108 4313
rect 5108 4264 5300 4304
rect 5068 4255 5108 4264
rect 4779 4220 4821 4229
rect 4779 4180 4780 4220
rect 4820 4180 4821 4220
rect 4779 4171 4821 4180
rect 4780 4136 4820 4171
rect 4780 4085 4820 4096
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 5067 4136 5109 4145
rect 5067 4096 5068 4136
rect 5108 4096 5109 4136
rect 5067 4087 5109 4096
rect 5260 4136 5300 4264
rect 5260 4087 5300 4096
rect 5644 4136 5684 4145
rect 5740 4136 5780 4768
rect 5932 4759 5972 4768
rect 5684 4096 5780 4136
rect 5644 4087 5684 4096
rect 4684 3928 4820 3968
rect 4587 3919 4629 3928
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4780 3632 4820 3928
rect 4492 3592 4820 3632
rect 4395 3548 4437 3557
rect 4395 3508 4396 3548
rect 4436 3508 4437 3548
rect 4395 3499 4437 3508
rect 4300 3464 4340 3473
rect 4204 3424 4300 3464
rect 4300 3415 4340 3424
rect 4396 3414 4436 3499
rect 4492 3464 4532 3592
rect 4876 3557 4916 4087
rect 5068 4002 5108 4087
rect 4875 3548 4917 3557
rect 4875 3508 4876 3548
rect 4916 3508 4917 3548
rect 4875 3499 4917 3508
rect 4492 3415 4532 3424
rect 2956 2836 3052 2876
rect 3052 2827 3092 2836
rect 3244 2836 3572 2876
rect 2804 2584 2900 2624
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 2764 2575 2804 2584
rect 3051 2575 3093 2584
rect 3244 2624 3284 2836
rect 6028 2633 6068 4936
rect 6316 4145 6356 5608
rect 6507 5060 6549 5069
rect 6507 5020 6508 5060
rect 6548 5020 6549 5060
rect 6507 5011 6549 5020
rect 6315 4136 6357 4145
rect 6315 4096 6316 4136
rect 6356 4096 6357 4136
rect 6315 4087 6357 4096
rect 6508 4136 6548 5011
rect 7660 4313 7700 8455
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 42988 8093 43028 9547
rect 43084 9353 43124 9631
rect 43083 9344 43125 9353
rect 43083 9304 43084 9344
rect 43124 9304 43125 9344
rect 43083 9295 43125 9304
rect 42987 8084 43029 8093
rect 42987 8044 42988 8084
rect 43028 8044 43029 8084
rect 42987 8035 43029 8044
rect 43276 7757 43316 9883
rect 43852 9521 43892 10060
rect 44427 10100 44469 10109
rect 44427 10060 44428 10100
rect 44468 10060 44469 10100
rect 44427 10051 44469 10060
rect 44428 9966 44468 10051
rect 44524 9521 44564 10144
rect 46252 10184 46292 10219
rect 46252 10133 46292 10144
rect 46444 10184 46484 10193
rect 46347 10100 46389 10109
rect 46347 10060 46348 10100
rect 46388 10060 46389 10100
rect 46347 10051 46389 10060
rect 46348 9966 46388 10051
rect 43851 9512 43893 9521
rect 43851 9472 43852 9512
rect 43892 9472 43893 9512
rect 43851 9463 43893 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 45867 9512 45909 9521
rect 45867 9472 45868 9512
rect 45908 9472 45909 9512
rect 45867 9463 45909 9472
rect 46060 9512 46100 9521
rect 43852 8924 43892 9463
rect 45387 9428 45429 9437
rect 45387 9388 45388 9428
rect 45428 9388 45429 9428
rect 45387 9379 45429 9388
rect 44716 9344 44756 9353
rect 44620 9304 44716 9344
rect 43948 8924 43988 8933
rect 43852 8884 43948 8924
rect 43948 8875 43988 8884
rect 44620 8672 44660 9304
rect 44716 9295 44756 9304
rect 44907 9260 44949 9269
rect 44907 9220 44908 9260
rect 44948 9220 44949 9260
rect 44907 9211 44949 9220
rect 44620 8623 44660 8632
rect 44236 8588 44276 8597
rect 43948 8504 43988 8513
rect 43988 8464 44180 8504
rect 43948 8455 43988 8464
rect 44140 8000 44180 8464
rect 44236 8177 44276 8548
rect 44235 8168 44277 8177
rect 44235 8128 44236 8168
rect 44276 8128 44277 8168
rect 44235 8119 44277 8128
rect 44428 8009 44468 8094
rect 44140 7951 44180 7960
rect 44236 8000 44276 8009
rect 44236 7757 44276 7960
rect 44427 8000 44469 8009
rect 44427 7960 44428 8000
rect 44468 7960 44469 8000
rect 44427 7951 44469 7960
rect 44812 8000 44852 8009
rect 44812 7841 44852 7960
rect 44908 8000 44948 9211
rect 45003 8168 45045 8177
rect 45003 8128 45004 8168
rect 45044 8128 45045 8168
rect 45388 8168 45428 9379
rect 45868 9378 45908 9463
rect 45579 9344 45621 9353
rect 45579 9304 45580 9344
rect 45620 9304 45621 9344
rect 46060 9344 46100 9472
rect 46252 9344 46292 9353
rect 46060 9304 46252 9344
rect 45579 9295 45621 9304
rect 46252 9295 46292 9304
rect 45483 8756 45525 8765
rect 45483 8716 45484 8756
rect 45524 8716 45525 8756
rect 45483 8707 45525 8716
rect 45484 8672 45524 8707
rect 45484 8621 45524 8632
rect 45388 8128 45524 8168
rect 45003 8119 45045 8128
rect 45004 8034 45044 8119
rect 44908 7951 44948 7960
rect 45100 8000 45140 8009
rect 45388 8000 45428 8009
rect 45140 7960 45388 8000
rect 45100 7951 45140 7960
rect 45388 7951 45428 7960
rect 45484 8000 45524 8128
rect 44427 7832 44469 7841
rect 44427 7792 44428 7832
rect 44468 7792 44469 7832
rect 44427 7783 44469 7792
rect 44811 7832 44853 7841
rect 44811 7792 44812 7832
rect 44852 7792 44853 7832
rect 44811 7783 44853 7792
rect 43275 7748 43317 7757
rect 43275 7708 43276 7748
rect 43316 7708 43317 7748
rect 43275 7699 43317 7708
rect 44235 7748 44277 7757
rect 44235 7708 44236 7748
rect 44276 7708 44277 7748
rect 44235 7699 44277 7708
rect 44428 7698 44468 7783
rect 45387 7748 45429 7757
rect 45387 7708 45388 7748
rect 45428 7708 45429 7748
rect 45387 7699 45429 7708
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 45388 7160 45428 7699
rect 45388 7111 45428 7120
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 45484 6413 45524 7960
rect 45580 8000 45620 9295
rect 46444 9269 46484 10144
rect 46540 10184 46580 10396
rect 46827 10387 46869 10396
rect 46540 10135 46580 10144
rect 46731 10100 46773 10109
rect 46731 10060 46732 10100
rect 46772 10060 46773 10100
rect 46731 10051 46773 10060
rect 46732 9966 46772 10051
rect 46540 9512 46580 9521
rect 45963 9260 46005 9269
rect 45963 9220 45964 9260
rect 46004 9220 46005 9260
rect 45963 9211 46005 9220
rect 46443 9260 46485 9269
rect 46443 9220 46444 9260
rect 46484 9220 46485 9260
rect 46443 9211 46485 9220
rect 45964 9126 46004 9211
rect 46540 8924 46580 9472
rect 46636 9512 46676 9521
rect 46828 9512 46868 10387
rect 46924 10184 46964 10984
rect 47116 11024 47156 11033
rect 47116 10445 47156 10984
rect 48076 10974 48116 11059
rect 48460 11024 48500 11033
rect 48172 10984 48460 11024
rect 47884 10856 47924 10865
rect 48172 10856 48212 10984
rect 48460 10975 48500 10984
rect 49323 11024 49365 11033
rect 49323 10984 49324 11024
rect 49364 10984 49365 11024
rect 49323 10975 49365 10984
rect 49324 10890 49364 10975
rect 47924 10816 48212 10856
rect 47884 10807 47924 10816
rect 47115 10436 47157 10445
rect 47115 10396 47116 10436
rect 47156 10396 47157 10436
rect 47115 10387 47157 10396
rect 49131 10436 49173 10445
rect 49131 10396 49132 10436
rect 49172 10396 49173 10436
rect 49131 10387 49173 10396
rect 48363 10352 48405 10361
rect 48363 10312 48364 10352
rect 48404 10312 48405 10352
rect 48363 10303 48405 10312
rect 47116 10184 47156 10193
rect 46924 10144 47060 10184
rect 46923 9932 46965 9941
rect 46923 9892 46924 9932
rect 46964 9892 46965 9932
rect 46923 9883 46965 9892
rect 46676 9472 46868 9512
rect 46924 9512 46964 9883
rect 46636 9463 46676 9472
rect 46636 8924 46676 8933
rect 46540 8884 46636 8924
rect 46636 8875 46676 8884
rect 46539 8756 46581 8765
rect 46539 8716 46540 8756
rect 46580 8716 46581 8756
rect 46539 8707 46581 8716
rect 45483 6404 45525 6413
rect 45483 6364 45484 6404
rect 45524 6364 45525 6404
rect 45483 6355 45525 6364
rect 45580 6329 45620 7960
rect 45675 8000 45717 8009
rect 45675 7960 45676 8000
rect 45716 7960 45717 8000
rect 45675 7951 45717 7960
rect 45676 7866 45716 7951
rect 45868 7832 45908 7841
rect 45772 7160 45812 7169
rect 45868 7160 45908 7792
rect 45812 7120 45908 7160
rect 46540 7160 46580 8707
rect 46924 8597 46964 9472
rect 46923 8588 46965 8597
rect 46923 8548 46924 8588
rect 46964 8548 46965 8588
rect 46923 8539 46965 8548
rect 46636 8504 46676 8513
rect 46676 8464 46772 8504
rect 46636 8455 46676 8464
rect 46732 8009 46772 8464
rect 47020 8420 47060 10144
rect 47116 9344 47156 10144
rect 47980 10184 48020 10195
rect 47212 9344 47252 9353
rect 47116 9304 47212 9344
rect 47212 9295 47252 9304
rect 47980 8765 48020 10144
rect 47979 8756 48021 8765
rect 47979 8716 47980 8756
rect 48020 8716 48021 8756
rect 47979 8707 48021 8716
rect 48171 8756 48213 8765
rect 48171 8716 48172 8756
rect 48212 8716 48213 8756
rect 48171 8707 48213 8716
rect 47979 8588 48021 8597
rect 47979 8548 47980 8588
rect 48020 8548 48021 8588
rect 47979 8539 48021 8548
rect 46828 8380 47060 8420
rect 46731 8000 46773 8009
rect 46731 7960 46732 8000
rect 46772 7960 46773 8000
rect 46731 7951 46773 7960
rect 46828 8000 46868 8380
rect 47020 8009 47060 8094
rect 46732 7866 46772 7951
rect 46828 7841 46868 7960
rect 47019 8000 47061 8009
rect 47019 7960 47020 8000
rect 47060 7960 47061 8000
rect 47019 7951 47061 7960
rect 47212 8000 47252 8009
rect 46827 7832 46869 7841
rect 46827 7792 46828 7832
rect 46868 7792 46869 7832
rect 46827 7783 46869 7792
rect 47020 7832 47060 7841
rect 47212 7832 47252 7960
rect 47307 8000 47349 8009
rect 47500 8000 47540 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 47404 7960 47500 8000
rect 47308 7866 47348 7951
rect 47060 7792 47252 7832
rect 47020 7783 47060 7792
rect 46636 7160 46676 7169
rect 46540 7120 46636 7160
rect 46676 7120 46964 7160
rect 45772 7111 45812 7120
rect 46636 7111 46676 7120
rect 45579 6320 45621 6329
rect 45579 6280 45580 6320
rect 45620 6280 45621 6320
rect 45579 6271 45621 6280
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 46156 5816 46196 5825
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 45675 5060 45717 5069
rect 45675 5020 45676 5060
rect 45716 5020 45717 5060
rect 45675 5011 45717 5020
rect 45676 4926 45716 5011
rect 46060 4976 46100 4985
rect 46156 4976 46196 5776
rect 46100 4936 46196 4976
rect 46924 4976 46964 7120
rect 47212 6656 47252 6665
rect 47404 6656 47444 7960
rect 47500 7951 47540 7960
rect 47980 8000 48020 8539
rect 48020 7960 48116 8000
rect 47980 7951 48020 7960
rect 47691 7916 47733 7925
rect 47691 7876 47692 7916
rect 47732 7876 47733 7916
rect 47691 7867 47733 7876
rect 47499 7748 47541 7757
rect 47499 7708 47500 7748
rect 47540 7708 47541 7748
rect 47499 7699 47541 7708
rect 47500 7614 47540 7699
rect 47499 7412 47541 7421
rect 47499 7372 47500 7412
rect 47540 7372 47541 7412
rect 47499 7363 47541 7372
rect 47252 6616 47444 6656
rect 47212 6607 47252 6616
rect 47308 6488 47348 6499
rect 47308 6413 47348 6448
rect 47404 6488 47444 6497
rect 47115 6404 47157 6413
rect 47115 6364 47116 6404
rect 47156 6364 47157 6404
rect 47115 6355 47157 6364
rect 47307 6404 47349 6413
rect 47307 6364 47308 6404
rect 47348 6364 47349 6404
rect 47307 6355 47349 6364
rect 46060 4927 46100 4936
rect 46924 4927 46964 4936
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 7659 4304 7701 4313
rect 7659 4264 7660 4304
rect 7700 4264 7701 4304
rect 7659 4255 7701 4264
rect 7660 4170 7700 4255
rect 6508 4087 6548 4096
rect 47116 3968 47156 6355
rect 47404 6329 47444 6448
rect 47500 6488 47540 7363
rect 47500 6439 47540 6448
rect 47692 6488 47732 7867
rect 47883 7832 47925 7841
rect 47883 7792 47884 7832
rect 47924 7792 47925 7832
rect 47883 7783 47925 7792
rect 47787 7412 47829 7421
rect 47787 7372 47788 7412
rect 47828 7372 47829 7412
rect 47787 7363 47829 7372
rect 47788 7278 47828 7363
rect 47692 6439 47732 6448
rect 47884 6488 47924 7783
rect 47979 7412 48021 7421
rect 47979 7372 47980 7412
rect 48020 7372 48021 7412
rect 47979 7363 48021 7372
rect 47403 6320 47445 6329
rect 47403 6280 47404 6320
rect 47444 6280 47445 6320
rect 47403 6271 47445 6280
rect 47404 5825 47444 6271
rect 47692 6236 47732 6245
rect 47500 6196 47692 6236
rect 47403 5816 47445 5825
rect 47403 5776 47404 5816
rect 47444 5776 47445 5816
rect 47403 5767 47445 5776
rect 47212 5648 47252 5657
rect 47212 4808 47252 5608
rect 47403 5648 47445 5657
rect 47403 5608 47404 5648
rect 47444 5608 47445 5648
rect 47403 5599 47445 5608
rect 47500 5648 47540 6196
rect 47692 6187 47732 6196
rect 47595 5816 47637 5825
rect 47595 5776 47596 5816
rect 47636 5776 47637 5816
rect 47595 5767 47637 5776
rect 47500 5599 47540 5608
rect 47404 5514 47444 5599
rect 47308 5480 47348 5489
rect 47308 5069 47348 5440
rect 47307 5060 47349 5069
rect 47307 5020 47308 5060
rect 47348 5020 47349 5060
rect 47307 5011 47349 5020
rect 47212 4768 47444 4808
rect 47404 4136 47444 4768
rect 47404 4087 47444 4096
rect 47500 4136 47540 4145
rect 47500 3968 47540 4096
rect 47596 4136 47636 5767
rect 47884 5489 47924 6448
rect 47980 6488 48020 7363
rect 47980 6439 48020 6448
rect 48076 5648 48116 7960
rect 48172 6488 48212 8707
rect 48364 8504 48404 10303
rect 49132 10302 49172 10387
rect 48843 10268 48885 10277
rect 48843 10228 48844 10268
rect 48884 10228 48885 10268
rect 48843 10219 48885 10228
rect 48459 9512 48501 9521
rect 48459 9472 48460 9512
rect 48500 9472 48501 9512
rect 48459 9463 48501 9472
rect 48460 8765 48500 9463
rect 48459 8756 48501 8765
rect 48459 8716 48460 8756
rect 48500 8716 48501 8756
rect 48459 8707 48501 8716
rect 48460 8672 48500 8707
rect 48460 8622 48500 8632
rect 48652 8672 48692 8681
rect 48555 8588 48597 8597
rect 48555 8548 48556 8588
rect 48596 8548 48597 8588
rect 48555 8539 48597 8548
rect 48364 8464 48500 8504
rect 48267 8252 48309 8261
rect 48267 8212 48268 8252
rect 48308 8212 48309 8252
rect 48267 8203 48309 8212
rect 48268 8000 48308 8203
rect 48268 7951 48308 7960
rect 48364 8000 48404 8009
rect 48364 7421 48404 7960
rect 48460 7664 48500 8464
rect 48556 8009 48596 8539
rect 48555 8000 48597 8009
rect 48555 7960 48556 8000
rect 48596 7960 48597 8000
rect 48555 7951 48597 7960
rect 48652 7832 48692 8632
rect 48844 8672 48884 10219
rect 49804 9344 49844 11479
rect 49996 11033 50036 15259
rect 50188 11780 50228 15688
rect 50284 11957 50324 16780
rect 50476 16745 50516 17779
rect 50475 16736 50517 16745
rect 50475 16696 50476 16736
rect 50516 16696 50517 16736
rect 50475 16687 50517 16696
rect 50379 15392 50421 15401
rect 50379 15352 50380 15392
rect 50420 15352 50421 15392
rect 50379 15343 50421 15352
rect 50380 14972 50420 15343
rect 50380 14923 50420 14932
rect 50572 14393 50612 17863
rect 50668 17744 50708 17753
rect 50764 17744 50804 18376
rect 50708 17704 50804 17744
rect 50668 17695 50708 17704
rect 50667 17240 50709 17249
rect 50667 17200 50668 17240
rect 50708 17200 50709 17240
rect 50667 17191 50709 17200
rect 50668 17072 50708 17191
rect 50668 17023 50708 17032
rect 50764 17072 50804 17081
rect 50764 15569 50804 17032
rect 50860 16661 50900 18787
rect 51340 18500 51380 18511
rect 51340 18425 51380 18460
rect 51339 18416 51381 18425
rect 51339 18376 51340 18416
rect 51380 18376 51381 18416
rect 51339 18367 51381 18376
rect 51148 18332 51188 18341
rect 51148 17072 51188 18292
rect 51340 17333 51380 18367
rect 51532 17744 51572 17753
rect 51339 17324 51381 17333
rect 51339 17284 51340 17324
rect 51380 17284 51381 17324
rect 51339 17275 51381 17284
rect 51435 17240 51477 17249
rect 51435 17200 51436 17240
rect 51476 17200 51477 17240
rect 51435 17191 51477 17200
rect 51339 17156 51381 17165
rect 51339 17116 51340 17156
rect 51380 17116 51381 17156
rect 51339 17107 51381 17116
rect 51244 17072 51284 17081
rect 50956 17032 51244 17072
rect 50859 16652 50901 16661
rect 50859 16612 50860 16652
rect 50900 16612 50901 16652
rect 50859 16603 50901 16612
rect 50763 15560 50805 15569
rect 50850 15567 50890 15576
rect 50763 15520 50764 15560
rect 50804 15527 50850 15560
rect 50804 15520 50890 15527
rect 50763 15511 50805 15520
rect 50850 15518 50890 15520
rect 50956 15560 50996 17032
rect 51244 17023 51284 17032
rect 51340 17022 51380 17107
rect 51436 17072 51476 17191
rect 51436 17023 51476 17032
rect 51339 16904 51381 16913
rect 51339 16864 51340 16904
rect 51380 16864 51381 16904
rect 51339 16855 51381 16864
rect 51052 16820 51092 16829
rect 51052 16232 51092 16780
rect 51340 16484 51380 16855
rect 51340 16435 51380 16444
rect 51244 16232 51284 16241
rect 51052 16192 51244 16232
rect 51244 16183 51284 16192
rect 51436 16232 51476 16241
rect 51532 16232 51572 17704
rect 51628 17001 51668 19963
rect 51723 18332 51765 18341
rect 51723 18292 51724 18332
rect 51764 18292 51765 18332
rect 51916 18332 51956 25087
rect 52012 24464 52052 25171
rect 52108 24977 52148 25264
rect 52204 25852 52588 25892
rect 52107 24968 52149 24977
rect 52107 24928 52108 24968
rect 52148 24928 52149 24968
rect 52107 24919 52149 24928
rect 52204 24800 52244 25852
rect 52588 25843 52628 25852
rect 52683 25892 52725 25901
rect 52683 25852 52684 25892
rect 52724 25852 52725 25892
rect 52683 25843 52725 25852
rect 52684 25313 52724 25843
rect 52683 25304 52725 25313
rect 52683 25264 52684 25304
rect 52724 25264 52725 25304
rect 52683 25255 52725 25264
rect 52780 25304 52820 25936
rect 52876 25927 52916 25936
rect 52875 25640 52917 25649
rect 52875 25600 52876 25640
rect 52916 25600 52917 25640
rect 52875 25591 52917 25600
rect 52780 25255 52820 25264
rect 52395 25220 52437 25229
rect 52395 25180 52396 25220
rect 52436 25180 52437 25220
rect 52395 25171 52437 25180
rect 52396 25086 52436 25171
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 52204 24760 52436 24800
rect 52108 24632 52148 24641
rect 52299 24632 52341 24641
rect 52148 24592 52244 24632
rect 52108 24583 52148 24592
rect 52204 24473 52244 24592
rect 52299 24592 52300 24632
rect 52340 24592 52341 24632
rect 52299 24583 52341 24592
rect 52396 24632 52436 24760
rect 52396 24583 52436 24592
rect 52300 24498 52340 24583
rect 52108 24464 52148 24473
rect 52012 24424 52108 24464
rect 52108 24415 52148 24424
rect 52203 24464 52245 24473
rect 52203 24424 52204 24464
rect 52244 24424 52245 24464
rect 52203 24415 52245 24424
rect 52588 24464 52628 24473
rect 52204 23969 52244 24415
rect 52203 23960 52245 23969
rect 52203 23920 52204 23960
rect 52244 23920 52245 23960
rect 52203 23911 52245 23920
rect 52108 23792 52148 23801
rect 52588 23792 52628 24424
rect 52148 23752 52628 23792
rect 52108 23743 52148 23752
rect 52876 23708 52916 25591
rect 53164 24473 53204 28111
rect 53292 27656 53334 27665
rect 53292 27616 53293 27656
rect 53333 27616 53334 27656
rect 53292 27607 53334 27616
rect 53293 27497 53333 27607
rect 53292 27488 53334 27497
rect 53292 27448 53293 27488
rect 53333 27448 53334 27488
rect 53292 27439 53334 27448
rect 54219 27068 54261 27077
rect 54219 27028 54220 27068
rect 54260 27028 54261 27068
rect 54219 27019 54261 27028
rect 54220 26934 54260 27019
rect 53644 25304 53684 25313
rect 53644 24641 53684 25264
rect 53643 24632 53685 24641
rect 53643 24592 53644 24632
rect 53684 24592 53685 24632
rect 53643 24583 53685 24592
rect 53163 24464 53205 24473
rect 53163 24424 53164 24464
rect 53204 24424 53205 24464
rect 53163 24415 53205 24424
rect 53644 23801 53684 24583
rect 54316 24557 54356 29623
rect 54699 28832 54741 28841
rect 54699 28792 54700 28832
rect 54740 28792 54741 28832
rect 54699 28783 54741 28792
rect 54603 28580 54645 28589
rect 54603 28540 54604 28580
rect 54644 28540 54645 28580
rect 54603 28531 54645 28540
rect 54507 28496 54549 28505
rect 54507 28456 54508 28496
rect 54548 28456 54549 28496
rect 54507 28447 54549 28456
rect 54508 27488 54548 28447
rect 54604 28446 54644 28531
rect 54604 27656 54644 27665
rect 54700 27656 54740 28783
rect 54892 28757 54932 30808
rect 54988 30269 55028 32320
rect 55179 32108 55221 32117
rect 55179 32068 55180 32108
rect 55220 32068 55221 32108
rect 55179 32059 55221 32068
rect 55180 31604 55220 32059
rect 55180 31555 55220 31564
rect 55372 31436 55412 33319
rect 55660 33209 55700 35428
rect 55948 35384 55988 35848
rect 56043 35888 56085 35897
rect 56043 35848 56044 35888
rect 56084 35848 56085 35888
rect 56043 35839 56085 35848
rect 56236 35888 56276 36595
rect 55756 35344 55988 35384
rect 55659 33200 55701 33209
rect 55659 33160 55660 33200
rect 55700 33160 55701 33200
rect 55659 33151 55701 33160
rect 55468 33032 55508 33041
rect 55508 32992 55700 33032
rect 55468 32983 55508 32992
rect 55468 32864 55508 32873
rect 55468 31445 55508 32824
rect 55660 32864 55700 32992
rect 55660 32815 55700 32824
rect 55563 32528 55605 32537
rect 55563 32488 55564 32528
rect 55604 32488 55605 32528
rect 55563 32479 55605 32488
rect 55084 31396 55412 31436
rect 55467 31436 55509 31445
rect 55467 31396 55468 31436
rect 55508 31396 55509 31436
rect 55084 30680 55124 31396
rect 55467 31387 55509 31396
rect 55564 31352 55604 32479
rect 55756 31949 55796 35344
rect 55948 35216 55988 35225
rect 55851 35132 55893 35141
rect 55851 35092 55852 35132
rect 55892 35092 55893 35132
rect 55851 35083 55893 35092
rect 55852 34376 55892 35083
rect 55948 34553 55988 35176
rect 56044 35141 56084 35839
rect 56043 35132 56085 35141
rect 56043 35092 56044 35132
rect 56084 35092 56085 35132
rect 56043 35083 56085 35092
rect 56236 34628 56276 35848
rect 56428 35888 56468 35897
rect 56331 35804 56373 35813
rect 56331 35764 56332 35804
rect 56372 35764 56373 35804
rect 56331 35755 56373 35764
rect 56332 35670 56372 35755
rect 56428 34889 56468 35848
rect 56619 35720 56661 35729
rect 56619 35680 56620 35720
rect 56660 35680 56661 35720
rect 56619 35671 56661 35680
rect 56620 35586 56660 35671
rect 56716 35216 56756 37183
rect 57099 36896 57141 36905
rect 57099 36856 57100 36896
rect 57140 36856 57141 36896
rect 57099 36847 57141 36856
rect 57100 36762 57140 36847
rect 57004 36728 57044 36737
rect 56812 36476 56852 36485
rect 56852 36436 56948 36476
rect 56812 36427 56852 36436
rect 56811 35972 56853 35981
rect 56811 35932 56812 35972
rect 56852 35932 56853 35972
rect 56811 35923 56853 35932
rect 56812 35838 56852 35923
rect 56908 35897 56948 36436
rect 56907 35888 56949 35897
rect 56907 35848 56908 35888
rect 56948 35848 56949 35888
rect 56907 35839 56949 35848
rect 57004 35225 57044 36688
rect 57196 36728 57236 36739
rect 57196 36653 57236 36688
rect 57291 36728 57333 36737
rect 57291 36688 57292 36728
rect 57332 36688 57333 36728
rect 57291 36679 57333 36688
rect 57195 36644 57237 36653
rect 57195 36604 57196 36644
rect 57236 36604 57237 36644
rect 57195 36595 57237 36604
rect 57292 36594 57332 36679
rect 56812 35216 56852 35225
rect 56716 35176 56812 35216
rect 56427 34880 56469 34889
rect 56427 34840 56428 34880
rect 56468 34840 56469 34880
rect 56427 34831 56469 34840
rect 56236 34588 56372 34628
rect 55947 34544 55989 34553
rect 55947 34504 55948 34544
rect 55988 34504 55989 34544
rect 55947 34495 55989 34504
rect 55852 34327 55892 34336
rect 55947 34376 55989 34385
rect 55947 34336 55948 34376
rect 55988 34336 55989 34376
rect 55947 34327 55989 34336
rect 56235 34376 56277 34385
rect 56235 34336 56236 34376
rect 56276 34336 56277 34376
rect 56235 34327 56277 34336
rect 55948 34242 55988 34327
rect 56236 34049 56276 34327
rect 56332 34301 56372 34588
rect 56428 34469 56468 34831
rect 56523 34544 56565 34553
rect 56523 34504 56524 34544
rect 56564 34504 56565 34544
rect 56523 34495 56565 34504
rect 56427 34460 56469 34469
rect 56427 34420 56428 34460
rect 56468 34420 56469 34460
rect 56427 34411 56469 34420
rect 56524 34410 56564 34495
rect 56331 34292 56373 34301
rect 56331 34252 56332 34292
rect 56372 34252 56373 34292
rect 56331 34243 56373 34252
rect 55851 34040 55893 34049
rect 55851 34000 55852 34040
rect 55892 34000 55893 34040
rect 55851 33991 55893 34000
rect 56235 34040 56277 34049
rect 56235 34000 56236 34040
rect 56276 34000 56277 34040
rect 56235 33991 56277 34000
rect 55852 33140 55892 33991
rect 56140 33536 56180 33545
rect 56140 33140 56180 33496
rect 56332 33293 56372 34243
rect 56331 33284 56373 33293
rect 56331 33244 56332 33284
rect 56372 33244 56373 33284
rect 56331 33235 56373 33244
rect 55852 33100 55988 33140
rect 55755 31940 55797 31949
rect 55755 31900 55756 31940
rect 55796 31900 55892 31940
rect 55755 31891 55797 31900
rect 55180 31184 55220 31193
rect 55220 31144 55508 31184
rect 55180 31135 55220 31144
rect 55275 31016 55317 31025
rect 55275 30976 55276 31016
rect 55316 30976 55317 31016
rect 55275 30967 55317 30976
rect 55084 30437 55124 30640
rect 55083 30428 55125 30437
rect 55083 30388 55084 30428
rect 55124 30388 55125 30428
rect 55083 30379 55125 30388
rect 54987 30260 55029 30269
rect 54987 30220 54988 30260
rect 55028 30220 55029 30260
rect 54987 30211 55029 30220
rect 55179 29924 55221 29933
rect 55179 29884 55180 29924
rect 55220 29884 55221 29924
rect 55179 29875 55221 29884
rect 54987 29840 55029 29849
rect 54987 29800 54988 29840
rect 55028 29800 55029 29840
rect 54987 29791 55029 29800
rect 55084 29840 55124 29849
rect 54988 29706 55028 29791
rect 54987 29588 55029 29597
rect 54987 29548 54988 29588
rect 55028 29548 55029 29588
rect 54987 29539 55029 29548
rect 54891 28748 54933 28757
rect 54891 28708 54892 28748
rect 54932 28708 54933 28748
rect 54891 28699 54933 28708
rect 54892 28253 54932 28699
rect 54891 28244 54933 28253
rect 54891 28204 54892 28244
rect 54932 28204 54933 28244
rect 54891 28195 54933 28204
rect 54644 27616 54740 27656
rect 54795 27656 54837 27665
rect 54795 27616 54796 27656
rect 54836 27616 54837 27656
rect 54604 27607 54644 27616
rect 54795 27607 54837 27616
rect 54892 27656 54932 27665
rect 54796 27522 54836 27607
rect 54604 27488 54644 27497
rect 54508 27448 54604 27488
rect 54604 27439 54644 27448
rect 54412 27404 54452 27413
rect 54412 26741 54452 27364
rect 54892 27329 54932 27616
rect 54891 27320 54933 27329
rect 54891 27280 54892 27320
rect 54932 27280 54933 27320
rect 54891 27271 54933 27280
rect 54411 26732 54453 26741
rect 54411 26692 54412 26732
rect 54452 26692 54453 26732
rect 54411 26683 54453 26692
rect 54699 26732 54741 26741
rect 54699 26692 54700 26732
rect 54740 26692 54741 26732
rect 54699 26683 54741 26692
rect 54700 26321 54740 26683
rect 54699 26312 54741 26321
rect 54699 26272 54700 26312
rect 54740 26272 54741 26312
rect 54699 26263 54741 26272
rect 54988 26144 55028 29539
rect 55084 29345 55124 29800
rect 55083 29336 55125 29345
rect 55083 29296 55084 29336
rect 55124 29296 55125 29336
rect 55083 29287 55125 29296
rect 55180 27656 55220 29875
rect 55276 29504 55316 30967
rect 55371 30764 55413 30773
rect 55371 30724 55372 30764
rect 55412 30724 55413 30764
rect 55371 30715 55413 30724
rect 55468 30764 55508 31144
rect 55468 30715 55508 30724
rect 55372 30680 55412 30715
rect 55372 30629 55412 30640
rect 55564 30260 55604 31312
rect 55756 31352 55796 31361
rect 55660 31268 55700 31277
rect 55660 30689 55700 31228
rect 55659 30680 55701 30689
rect 55659 30640 55660 30680
rect 55700 30640 55701 30680
rect 55659 30631 55701 30640
rect 55756 30512 55796 31312
rect 55756 30463 55796 30472
rect 55468 30220 55604 30260
rect 55468 29597 55508 30220
rect 55852 30176 55892 31900
rect 55948 31025 55988 33100
rect 56044 33100 56180 33140
rect 56332 33140 56372 33235
rect 56812 33140 56852 35176
rect 57003 35216 57045 35225
rect 57003 35176 57004 35216
rect 57044 35176 57045 35216
rect 57003 35167 57045 35176
rect 56332 33100 56468 33140
rect 56812 33100 56948 33140
rect 56044 32864 56084 33100
rect 56044 32815 56084 32824
rect 56140 31268 56180 31277
rect 55947 31016 55989 31025
rect 55947 30976 55948 31016
rect 55988 30976 55989 31016
rect 55947 30967 55989 30976
rect 55947 30848 55989 30857
rect 55947 30808 55948 30848
rect 55988 30808 55989 30848
rect 55947 30799 55989 30808
rect 56044 30848 56084 30857
rect 56140 30848 56180 31228
rect 56084 30808 56180 30848
rect 56044 30799 56084 30808
rect 55948 30680 55988 30799
rect 55948 30353 55988 30640
rect 56139 30680 56181 30689
rect 56139 30640 56140 30680
rect 56180 30640 56181 30680
rect 56139 30631 56181 30640
rect 56236 30680 56276 30691
rect 56140 30546 56180 30631
rect 56236 30605 56276 30640
rect 56428 30680 56468 33100
rect 56908 32864 56948 33100
rect 56620 32024 56660 32033
rect 56524 31984 56620 32024
rect 56524 31352 56564 31984
rect 56620 31975 56660 31984
rect 56908 31361 56948 32824
rect 56524 31303 56564 31312
rect 56907 31352 56949 31361
rect 56907 31312 56908 31352
rect 56948 31312 56949 31352
rect 56907 31303 56949 31312
rect 56619 31100 56661 31109
rect 56619 31060 56620 31100
rect 56660 31060 56661 31100
rect 56619 31051 56661 31060
rect 56620 30773 56660 31051
rect 56619 30764 56661 30773
rect 56619 30724 56620 30764
rect 56660 30724 56661 30764
rect 56619 30715 56661 30724
rect 56235 30596 56277 30605
rect 56235 30556 56236 30596
rect 56276 30556 56277 30596
rect 56235 30547 56277 30556
rect 55947 30344 55989 30353
rect 55947 30304 55948 30344
rect 55988 30304 55989 30344
rect 55947 30295 55989 30304
rect 56331 30344 56373 30353
rect 56331 30304 56332 30344
rect 56372 30304 56373 30344
rect 56331 30295 56373 30304
rect 56235 30260 56277 30269
rect 56235 30220 56236 30260
rect 56276 30220 56277 30260
rect 56235 30211 56277 30220
rect 55564 30136 55892 30176
rect 55467 29588 55509 29597
rect 55467 29548 55468 29588
rect 55508 29548 55509 29588
rect 55467 29539 55509 29548
rect 55276 29464 55412 29504
rect 55275 29336 55317 29345
rect 55275 29296 55276 29336
rect 55316 29296 55317 29336
rect 55275 29287 55317 29296
rect 55276 29202 55316 29287
rect 55275 28664 55317 28673
rect 55275 28624 55276 28664
rect 55316 28624 55317 28664
rect 55275 28615 55317 28624
rect 55180 27581 55220 27616
rect 55276 27656 55316 28615
rect 55372 28328 55412 29464
rect 55564 29420 55604 30136
rect 55756 30008 55796 30017
rect 55796 29968 55988 30008
rect 55756 29959 55796 29968
rect 55660 29840 55700 29849
rect 55660 29597 55700 29800
rect 55852 29840 55892 29849
rect 55659 29588 55701 29597
rect 55659 29548 55660 29588
rect 55700 29548 55701 29588
rect 55659 29539 55701 29548
rect 55564 29380 55700 29420
rect 55468 29168 55508 29177
rect 55468 28841 55508 29128
rect 55564 29168 55604 29177
rect 55467 28832 55509 28841
rect 55467 28792 55468 28832
rect 55508 28792 55509 28832
rect 55467 28783 55509 28792
rect 55564 28757 55604 29128
rect 55660 29168 55700 29380
rect 55755 29336 55797 29345
rect 55755 29296 55756 29336
rect 55796 29296 55797 29336
rect 55755 29287 55797 29296
rect 55563 28748 55605 28757
rect 55563 28708 55564 28748
rect 55604 28708 55605 28748
rect 55563 28699 55605 28708
rect 55564 28580 55604 28699
rect 55372 28169 55412 28288
rect 55468 28540 55604 28580
rect 55371 28160 55413 28169
rect 55371 28120 55372 28160
rect 55412 28120 55413 28160
rect 55371 28111 55413 28120
rect 55468 27917 55508 28540
rect 55660 28496 55700 29128
rect 55564 28456 55700 28496
rect 55756 29168 55796 29287
rect 55467 27908 55509 27917
rect 55467 27868 55468 27908
rect 55508 27868 55509 27908
rect 55467 27859 55509 27868
rect 55564 27824 55604 28456
rect 55659 28328 55701 28337
rect 55659 28288 55660 28328
rect 55700 28288 55701 28328
rect 55659 28279 55701 28288
rect 55756 28328 55796 29128
rect 55852 28580 55892 29800
rect 55948 28757 55988 29968
rect 56236 29924 56276 30211
rect 56236 29875 56276 29884
rect 56140 29168 56180 29177
rect 55947 28748 55989 28757
rect 55947 28708 55948 28748
rect 55988 28708 55989 28748
rect 55947 28699 55989 28708
rect 56044 28580 56084 28589
rect 55852 28540 56044 28580
rect 56140 28580 56180 29128
rect 56236 28580 56276 28589
rect 56140 28540 56236 28580
rect 56044 28531 56084 28540
rect 56236 28531 56276 28540
rect 55756 28279 55796 28288
rect 56236 28328 56276 28337
rect 56332 28328 56372 30295
rect 56428 30092 56468 30640
rect 56620 30680 56660 30715
rect 56620 30630 56660 30640
rect 56523 30596 56565 30605
rect 56523 30556 56524 30596
rect 56564 30556 56565 30596
rect 56523 30547 56565 30556
rect 56524 30462 56564 30547
rect 56428 29849 56468 30052
rect 56620 30008 56660 30017
rect 56427 29840 56469 29849
rect 56427 29800 56428 29840
rect 56468 29800 56469 29840
rect 56427 29791 56469 29800
rect 56524 29168 56564 29177
rect 56620 29168 56660 29968
rect 57004 29933 57044 35167
rect 57483 34964 57525 34973
rect 57483 34924 57484 34964
rect 57524 34924 57525 34964
rect 57483 34915 57525 34924
rect 57484 34376 57524 34915
rect 57484 34327 57524 34336
rect 57580 34376 57620 34385
rect 57580 33797 57620 34336
rect 57579 33788 57621 33797
rect 57579 33748 57580 33788
rect 57620 33748 57621 33788
rect 57579 33739 57621 33748
rect 57676 33041 57716 38116
rect 57867 38156 57909 38165
rect 57867 38116 57868 38156
rect 57908 38116 57909 38156
rect 57867 38107 57909 38116
rect 57868 38072 57908 38107
rect 57868 38021 57908 38032
rect 58059 37988 58101 37997
rect 58059 37948 58060 37988
rect 58100 37948 58101 37988
rect 58059 37939 58101 37948
rect 58060 37854 58100 37939
rect 58059 37316 58101 37325
rect 58059 37276 58060 37316
rect 58100 37276 58101 37316
rect 58059 37267 58101 37276
rect 57964 34964 58004 34975
rect 57964 34889 58004 34924
rect 57963 34880 58005 34889
rect 57963 34840 57964 34880
rect 58004 34840 58005 34880
rect 57963 34831 58005 34840
rect 57772 34544 57812 34553
rect 57812 34504 58004 34544
rect 57772 34495 57812 34504
rect 57772 34376 57812 34385
rect 57772 33965 57812 34336
rect 57964 34376 58004 34504
rect 57964 34327 58004 34336
rect 58060 34217 58100 37267
rect 58156 37241 58196 38200
rect 58155 37232 58197 37241
rect 58155 37192 58156 37232
rect 58196 37192 58197 37232
rect 58155 37183 58197 37192
rect 58252 36905 58292 38200
rect 58348 38240 58388 38249
rect 58348 37493 58388 38200
rect 59403 38240 59445 38249
rect 59403 38200 59404 38240
rect 59444 38200 59445 38240
rect 59403 38191 59445 38200
rect 63532 38240 63572 38249
rect 63724 38240 63764 38249
rect 63572 38200 63668 38240
rect 63532 38191 63572 38200
rect 59404 38106 59444 38191
rect 59980 38156 60020 38167
rect 59980 38081 60020 38116
rect 59979 38072 60021 38081
rect 59979 38032 59980 38072
rect 60020 38032 60021 38072
rect 59979 38023 60021 38032
rect 60172 38072 60212 38081
rect 58828 37988 58868 37997
rect 58347 37484 58389 37493
rect 58347 37444 58348 37484
rect 58388 37444 58389 37484
rect 58347 37435 58389 37444
rect 58540 37400 58580 37409
rect 58348 37232 58388 37241
rect 58540 37232 58580 37360
rect 58388 37192 58580 37232
rect 58636 37400 58676 37409
rect 58251 36896 58293 36905
rect 58251 36856 58252 36896
rect 58292 36856 58293 36896
rect 58251 36847 58293 36856
rect 58348 36737 58388 37192
rect 58539 36980 58581 36989
rect 58539 36940 58540 36980
rect 58580 36940 58581 36980
rect 58539 36931 58581 36940
rect 58252 36728 58292 36737
rect 58155 35216 58197 35225
rect 58155 35176 58156 35216
rect 58196 35176 58197 35216
rect 58155 35167 58197 35176
rect 58156 35082 58196 35167
rect 58155 34964 58197 34973
rect 58155 34924 58156 34964
rect 58196 34924 58197 34964
rect 58155 34915 58197 34924
rect 58156 34830 58196 34915
rect 58155 34628 58197 34637
rect 58155 34588 58156 34628
rect 58196 34588 58197 34628
rect 58155 34579 58197 34588
rect 58059 34208 58101 34217
rect 58059 34168 58060 34208
rect 58100 34168 58101 34208
rect 58059 34159 58101 34168
rect 57771 33956 57813 33965
rect 57771 33916 57772 33956
rect 57812 33916 57813 33956
rect 57771 33907 57813 33916
rect 57771 33788 57813 33797
rect 57771 33748 57772 33788
rect 57812 33748 57813 33788
rect 57771 33739 57813 33748
rect 57675 33032 57717 33041
rect 57675 32992 57676 33032
rect 57716 32992 57717 33032
rect 57675 32983 57717 32992
rect 57772 32873 57812 33739
rect 57771 32864 57813 32873
rect 57771 32824 57772 32864
rect 57812 32824 57813 32864
rect 57771 32815 57813 32824
rect 58156 32864 58196 34579
rect 58252 34385 58292 36688
rect 58347 36728 58389 36737
rect 58347 36688 58348 36728
rect 58388 36688 58389 36728
rect 58347 36679 58389 36688
rect 58540 36728 58580 36931
rect 58636 36896 58676 37360
rect 58732 37400 58772 37411
rect 58828 37409 58868 37948
rect 59787 37988 59829 37997
rect 59787 37948 59788 37988
rect 59828 37948 59829 37988
rect 59787 37939 59829 37948
rect 59788 37854 59828 37939
rect 58732 37325 58772 37360
rect 58827 37400 58869 37409
rect 58827 37360 58828 37400
rect 58868 37360 58869 37400
rect 58827 37351 58869 37360
rect 59500 37400 59540 37409
rect 60172 37400 60212 38032
rect 60459 38072 60501 38081
rect 60459 38032 60460 38072
rect 60500 38032 60501 38072
rect 60459 38023 60501 38032
rect 61900 38072 61940 38081
rect 60267 37484 60309 37493
rect 60267 37444 60268 37484
rect 60308 37444 60309 37484
rect 60267 37435 60309 37444
rect 59540 37360 60212 37400
rect 59500 37351 59540 37360
rect 58731 37316 58773 37325
rect 58731 37276 58732 37316
rect 58772 37276 58773 37316
rect 58731 37267 58773 37276
rect 59116 37316 59156 37325
rect 58827 37232 58869 37241
rect 58827 37192 58828 37232
rect 58868 37192 58869 37232
rect 58827 37183 58869 37192
rect 58828 37098 58868 37183
rect 59019 36896 59061 36905
rect 58636 36856 58772 36896
rect 58540 36679 58580 36688
rect 58635 36728 58677 36737
rect 58635 36688 58636 36728
rect 58676 36688 58677 36728
rect 58635 36679 58677 36688
rect 58636 36594 58676 36679
rect 58732 35897 58772 36856
rect 59019 36856 59020 36896
rect 59060 36856 59061 36896
rect 59116 36896 59156 37276
rect 59787 36980 59829 36989
rect 59787 36940 59788 36980
rect 59828 36940 59829 36980
rect 59787 36931 59829 36940
rect 59212 36896 59252 36905
rect 59116 36856 59212 36896
rect 59019 36847 59061 36856
rect 59212 36847 59252 36856
rect 59307 36896 59349 36905
rect 59307 36856 59308 36896
rect 59348 36856 59349 36896
rect 59307 36847 59349 36856
rect 59404 36856 59732 36896
rect 58924 36476 58964 36485
rect 58828 36436 58924 36476
rect 58443 35888 58485 35897
rect 58443 35848 58444 35888
rect 58484 35848 58485 35888
rect 58443 35839 58485 35848
rect 58731 35888 58773 35897
rect 58731 35848 58732 35888
rect 58772 35848 58773 35888
rect 58731 35839 58773 35848
rect 58828 35888 58868 36436
rect 58924 36427 58964 36436
rect 59020 36308 59060 36847
rect 58924 36268 59060 36308
rect 59116 36728 59156 36737
rect 58924 35972 58964 36268
rect 58924 35923 58964 35932
rect 58828 35839 58868 35848
rect 59020 35888 59060 35897
rect 58348 35216 58388 35225
rect 58348 34553 58388 35176
rect 58444 35216 58484 35839
rect 58444 35167 58484 35176
rect 58636 35048 58676 35057
rect 58347 34544 58389 34553
rect 58347 34504 58348 34544
rect 58388 34504 58389 34544
rect 58347 34495 58389 34504
rect 58251 34376 58293 34385
rect 58251 34336 58252 34376
rect 58292 34336 58293 34376
rect 58251 34327 58293 34336
rect 58348 34376 58388 34385
rect 58636 34376 58676 35008
rect 58388 34336 58676 34376
rect 58348 34327 58388 34336
rect 58732 34292 58772 35839
rect 58540 34252 58772 34292
rect 58827 34292 58869 34301
rect 58827 34252 58828 34292
rect 58868 34252 58869 34292
rect 58443 34208 58485 34217
rect 58443 34168 58444 34208
rect 58484 34168 58485 34208
rect 58443 34159 58485 34168
rect 58347 33956 58389 33965
rect 58347 33916 58348 33956
rect 58388 33916 58389 33956
rect 58347 33907 58389 33916
rect 58348 33872 58388 33907
rect 58348 33821 58388 33832
rect 58444 33704 58484 34159
rect 58444 33655 58484 33664
rect 58540 33704 58580 34252
rect 58827 34243 58869 34252
rect 58828 33704 58868 34243
rect 59020 33872 59060 35848
rect 59116 34637 59156 36688
rect 59308 36728 59348 36847
rect 59308 36679 59348 36688
rect 59404 36728 59444 36856
rect 59692 36812 59732 36856
rect 59692 36763 59732 36772
rect 59404 36679 59444 36688
rect 59596 36728 59636 36737
rect 59115 34628 59157 34637
rect 59115 34588 59116 34628
rect 59156 34588 59157 34628
rect 59115 34579 59157 34588
rect 59596 34469 59636 36688
rect 59788 36728 59828 36931
rect 60268 36896 60308 37435
rect 60363 37400 60405 37409
rect 60363 37360 60364 37400
rect 60404 37360 60405 37400
rect 60363 37351 60405 37360
rect 60364 37266 60404 37351
rect 60460 36896 60500 38023
rect 61131 37988 61173 37997
rect 61131 37948 61132 37988
rect 61172 37948 61173 37988
rect 61131 37939 61173 37948
rect 60460 36856 60596 36896
rect 60268 36847 60308 36856
rect 60172 36728 60212 36737
rect 59788 36679 59828 36688
rect 59884 36688 60172 36728
rect 59788 35216 59828 35225
rect 59788 34553 59828 35176
rect 59787 34544 59829 34553
rect 59787 34504 59788 34544
rect 59828 34504 59829 34544
rect 59787 34495 59829 34504
rect 59595 34460 59637 34469
rect 59595 34420 59596 34460
rect 59636 34420 59637 34460
rect 59595 34411 59637 34420
rect 59211 34376 59253 34385
rect 59211 34336 59212 34376
rect 59252 34336 59253 34376
rect 59211 34327 59253 34336
rect 59212 34242 59252 34327
rect 59020 33832 59156 33872
rect 58540 33655 58580 33664
rect 58636 33659 58676 33668
rect 58828 33655 58868 33664
rect 59020 33704 59060 33713
rect 58539 33452 58581 33461
rect 58539 33412 58540 33452
rect 58580 33412 58581 33452
rect 58539 33403 58581 33412
rect 58444 32873 58484 32958
rect 58252 32864 58292 32873
rect 58156 32824 58252 32864
rect 58060 32696 58100 32707
rect 58060 32621 58100 32656
rect 58059 32612 58101 32621
rect 58059 32572 58060 32612
rect 58100 32572 58101 32612
rect 58059 32563 58101 32572
rect 57387 31352 57429 31361
rect 57387 31312 57388 31352
rect 57428 31312 57429 31352
rect 57387 31303 57429 31312
rect 57388 31218 57428 31303
rect 58156 30857 58196 32824
rect 58252 32815 58292 32824
rect 58443 32864 58485 32873
rect 58443 32824 58444 32864
rect 58484 32824 58485 32864
rect 58443 32815 58485 32824
rect 58540 32864 58580 33403
rect 58636 33284 58676 33619
rect 58923 33452 58965 33461
rect 58923 33412 58924 33452
rect 58964 33412 58965 33452
rect 58923 33403 58965 33412
rect 58924 33318 58964 33403
rect 58731 33284 58773 33293
rect 58636 33244 58732 33284
rect 58772 33244 58773 33284
rect 58731 33235 58773 33244
rect 58732 33140 58772 33235
rect 58732 33100 58868 33140
rect 58540 32815 58580 32824
rect 58347 32780 58389 32789
rect 58347 32740 58348 32780
rect 58388 32740 58389 32780
rect 58347 32731 58389 32740
rect 58348 32646 58388 32731
rect 58347 32276 58389 32285
rect 58347 32236 58348 32276
rect 58388 32236 58389 32276
rect 58347 32227 58389 32236
rect 58348 32192 58388 32227
rect 58155 30848 58197 30857
rect 58155 30808 58156 30848
rect 58196 30808 58197 30848
rect 58155 30799 58197 30808
rect 57771 30764 57813 30773
rect 57771 30724 57772 30764
rect 57812 30724 57813 30764
rect 57771 30715 57813 30724
rect 57772 30630 57812 30715
rect 58156 30680 58196 30689
rect 58196 30640 58292 30680
rect 58156 30631 58196 30640
rect 58252 30008 58292 30640
rect 58348 30101 58388 32152
rect 58444 32117 58484 32815
rect 58731 32780 58773 32789
rect 58731 32740 58732 32780
rect 58772 32740 58773 32780
rect 58731 32731 58773 32740
rect 58732 32646 58772 32731
rect 58635 32528 58677 32537
rect 58828 32528 58868 33100
rect 59020 32537 59060 33664
rect 59116 33125 59156 33832
rect 59691 33704 59733 33713
rect 59691 33664 59692 33704
rect 59732 33664 59733 33704
rect 59691 33655 59733 33664
rect 59212 33536 59252 33545
rect 59115 33116 59157 33125
rect 59115 33076 59116 33116
rect 59156 33076 59157 33116
rect 59115 33067 59157 33076
rect 59116 32864 59156 32873
rect 59212 32864 59252 33496
rect 59403 33116 59445 33125
rect 59403 33076 59404 33116
rect 59444 33076 59445 33116
rect 59403 33067 59445 33076
rect 59156 32824 59252 32864
rect 59116 32815 59156 32824
rect 58635 32488 58636 32528
rect 58676 32488 58677 32528
rect 58635 32479 58677 32488
rect 58732 32488 58868 32528
rect 58636 32192 58676 32479
rect 58732 32276 58772 32488
rect 58828 32369 58868 32488
rect 59019 32528 59061 32537
rect 59019 32488 59020 32528
rect 59060 32488 59061 32528
rect 59019 32479 59061 32488
rect 58827 32360 58869 32369
rect 58827 32320 58828 32360
rect 58868 32320 58869 32360
rect 58827 32311 58869 32320
rect 58732 32227 58772 32236
rect 58443 32108 58485 32117
rect 58443 32068 58444 32108
rect 58484 32068 58485 32108
rect 58443 32059 58485 32068
rect 58636 31865 58676 32152
rect 59212 32192 59252 32201
rect 59020 32024 59060 32033
rect 59212 32024 59252 32152
rect 59404 32192 59444 33067
rect 59595 32360 59637 32369
rect 59595 32320 59596 32360
rect 59636 32320 59637 32360
rect 59595 32311 59637 32320
rect 59404 32143 59444 32152
rect 59596 32192 59636 32311
rect 59596 32143 59636 32152
rect 59692 32192 59732 33655
rect 59884 32192 59924 36688
rect 60172 36679 60212 36688
rect 60364 36728 60404 36737
rect 60268 36056 60308 36065
rect 60172 36016 60268 36056
rect 60172 35216 60212 36016
rect 60268 36007 60308 36016
rect 60364 35981 60404 36688
rect 60459 36728 60501 36737
rect 60459 36688 60460 36728
rect 60500 36688 60501 36728
rect 60459 36679 60501 36688
rect 60460 36594 60500 36679
rect 60556 36476 60596 36856
rect 60460 36436 60596 36476
rect 60363 35972 60405 35981
rect 60363 35932 60364 35972
rect 60404 35932 60405 35972
rect 60363 35923 60405 35932
rect 60172 35167 60212 35176
rect 60171 34460 60213 34469
rect 60171 34420 60172 34460
rect 60212 34420 60213 34460
rect 60171 34411 60213 34420
rect 59979 34376 60021 34385
rect 59979 34336 59980 34376
rect 60020 34336 60021 34376
rect 59979 34327 60021 34336
rect 59307 32108 59349 32117
rect 59307 32068 59308 32108
rect 59348 32068 59349 32108
rect 59307 32059 59349 32068
rect 59060 31984 59252 32024
rect 59020 31975 59060 31984
rect 59308 31974 59348 32059
rect 58635 31856 58677 31865
rect 58635 31816 58636 31856
rect 58676 31816 58677 31856
rect 58635 31807 58677 31816
rect 59115 31772 59157 31781
rect 59115 31732 59116 31772
rect 59156 31732 59157 31772
rect 59115 31723 59157 31732
rect 59019 31688 59061 31697
rect 59019 31648 59020 31688
rect 59060 31648 59061 31688
rect 59019 31639 59061 31648
rect 59020 31361 59060 31639
rect 59019 31352 59061 31361
rect 59019 31312 59020 31352
rect 59060 31312 59061 31352
rect 59019 31303 59061 31312
rect 58540 31184 58580 31195
rect 58540 31109 58580 31144
rect 58539 31100 58581 31109
rect 58539 31060 58540 31100
rect 58580 31060 58581 31100
rect 58539 31051 58581 31060
rect 59020 30691 59060 31303
rect 59020 30642 59060 30651
rect 58347 30092 58389 30101
rect 58347 30052 58348 30092
rect 58388 30052 58389 30092
rect 58347 30043 58389 30052
rect 58827 30092 58869 30101
rect 58827 30052 58828 30092
rect 58868 30052 58869 30092
rect 58827 30043 58869 30052
rect 58252 29959 58292 29968
rect 57003 29924 57045 29933
rect 57003 29884 57004 29924
rect 57044 29884 57045 29924
rect 57003 29875 57045 29884
rect 58828 29849 58868 30043
rect 59020 29911 59060 29920
rect 56715 29840 56757 29849
rect 56715 29800 56716 29840
rect 56756 29800 56757 29840
rect 56715 29791 56757 29800
rect 58827 29840 58869 29849
rect 58827 29800 58828 29840
rect 58868 29800 58869 29840
rect 58827 29791 58869 29800
rect 56564 29128 56660 29168
rect 56524 29119 56564 29128
rect 56427 28748 56469 28757
rect 56427 28708 56428 28748
rect 56468 28708 56469 28748
rect 56427 28699 56469 28708
rect 56276 28288 56372 28328
rect 56428 28328 56468 28699
rect 56236 28279 56276 28288
rect 55660 28194 55700 28279
rect 56043 28160 56085 28169
rect 56043 28120 56044 28160
rect 56084 28120 56085 28160
rect 56043 28111 56085 28120
rect 55851 27908 55893 27917
rect 55851 27868 55852 27908
rect 55892 27868 55893 27908
rect 55851 27859 55893 27868
rect 55564 27784 55796 27824
rect 55372 27656 55412 27665
rect 55276 27616 55372 27656
rect 55179 27572 55221 27581
rect 55179 27532 55180 27572
rect 55220 27532 55221 27572
rect 55179 27523 55221 27532
rect 55180 27404 55220 27413
rect 55180 27329 55220 27364
rect 55180 27320 55222 27329
rect 55180 27280 55181 27320
rect 55221 27280 55222 27320
rect 55180 27271 55222 27280
rect 54988 26069 55028 26104
rect 55180 26144 55220 26153
rect 54987 26060 55029 26069
rect 54987 26020 54988 26060
rect 55028 26020 55029 26060
rect 54987 26011 55029 26020
rect 55083 25976 55125 25985
rect 55083 25936 55084 25976
rect 55124 25936 55125 25976
rect 55180 25976 55220 26104
rect 55276 26121 55316 27616
rect 55372 27607 55412 27616
rect 55468 27656 55508 27665
rect 55660 27656 55700 27665
rect 55508 27616 55660 27656
rect 55371 27488 55413 27497
rect 55371 27448 55372 27488
rect 55412 27448 55413 27488
rect 55371 27439 55413 27448
rect 55372 26816 55412 27439
rect 55468 27077 55508 27616
rect 55660 27607 55700 27616
rect 55756 27656 55796 27784
rect 55467 27068 55509 27077
rect 55467 27028 55468 27068
rect 55508 27028 55509 27068
rect 55467 27019 55509 27028
rect 55659 27068 55701 27077
rect 55659 27028 55660 27068
rect 55700 27028 55701 27068
rect 55659 27019 55701 27028
rect 55372 26767 55412 26776
rect 55563 26648 55605 26657
rect 55563 26608 55564 26648
rect 55604 26608 55605 26648
rect 55563 26599 55605 26608
rect 55564 26153 55604 26599
rect 55660 26228 55700 27019
rect 55756 26993 55796 27616
rect 55852 27656 55892 27859
rect 55852 27607 55892 27616
rect 55948 27656 55988 27665
rect 55755 26984 55797 26993
rect 55755 26944 55756 26984
rect 55796 26944 55797 26984
rect 55755 26935 55797 26944
rect 55948 26825 55988 27616
rect 55947 26816 55989 26825
rect 55947 26776 55948 26816
rect 55988 26776 55989 26816
rect 55947 26767 55989 26776
rect 56044 26405 56084 28111
rect 56428 27665 56468 28288
rect 56524 28328 56564 28337
rect 56524 28160 56564 28288
rect 56716 28328 56756 29791
rect 57579 29504 57621 29513
rect 57579 29464 57580 29504
rect 57620 29464 57621 29504
rect 57579 29455 57621 29464
rect 57195 29420 57237 29429
rect 57195 29380 57196 29420
rect 57236 29380 57237 29420
rect 57195 29371 57237 29380
rect 56907 28664 56949 28673
rect 56907 28624 56908 28664
rect 56948 28624 56949 28664
rect 56907 28615 56949 28624
rect 56908 28337 56948 28615
rect 56716 28279 56756 28288
rect 56907 28328 56949 28337
rect 56907 28288 56908 28328
rect 56948 28288 56949 28328
rect 56907 28279 56949 28288
rect 56812 28244 56852 28253
rect 56812 28160 56852 28204
rect 56908 28194 56948 28279
rect 56524 28120 56852 28160
rect 56427 27656 56469 27665
rect 56427 27616 56428 27656
rect 56468 27616 56469 27656
rect 56427 27607 56469 27616
rect 56811 27572 56853 27581
rect 56811 27532 56812 27572
rect 56852 27532 56853 27572
rect 56811 27523 56853 27532
rect 56140 27488 56180 27497
rect 56180 27448 56276 27488
rect 56140 27439 56180 27448
rect 56236 26816 56276 27448
rect 56236 26767 56276 26776
rect 56331 26816 56373 26825
rect 56331 26776 56332 26816
rect 56372 26776 56373 26816
rect 56331 26767 56373 26776
rect 56043 26396 56085 26405
rect 56043 26356 56044 26396
rect 56084 26356 56085 26396
rect 56043 26347 56085 26356
rect 55660 26179 55700 26188
rect 55563 26144 55605 26153
rect 55276 26081 55499 26121
rect 55563 26104 55564 26144
rect 55604 26104 55605 26144
rect 55563 26095 55605 26104
rect 55756 26144 55796 26153
rect 56044 26144 56084 26347
rect 55796 26104 55988 26144
rect 55756 26095 55796 26104
rect 55372 25976 55412 25985
rect 55180 25936 55372 25976
rect 55459 25976 55499 26081
rect 55659 25976 55701 25985
rect 55459 25936 55508 25976
rect 55083 25927 55125 25936
rect 55372 25927 55412 25936
rect 54795 25892 54837 25901
rect 54795 25852 54796 25892
rect 54836 25852 54837 25892
rect 54795 25843 54837 25852
rect 54796 25556 54836 25843
rect 55084 25842 55124 25927
rect 54796 25507 54836 25516
rect 55468 25313 55508 25936
rect 55659 25936 55660 25976
rect 55700 25936 55701 25976
rect 55659 25927 55701 25936
rect 55564 25472 55604 25481
rect 55467 25304 55509 25313
rect 55467 25264 55468 25304
rect 55508 25264 55509 25304
rect 55467 25255 55509 25264
rect 54796 25136 54836 25145
rect 54796 24977 54836 25096
rect 54795 24968 54837 24977
rect 54795 24928 54796 24968
rect 54836 24928 54837 24968
rect 54795 24919 54837 24928
rect 55084 24632 55124 24641
rect 55468 24632 55508 24641
rect 55564 24632 55604 25432
rect 55124 24592 55412 24632
rect 55084 24583 55124 24592
rect 54315 24548 54357 24557
rect 54315 24508 54316 24548
rect 54356 24508 54357 24548
rect 54315 24499 54357 24508
rect 55275 24464 55317 24473
rect 55275 24424 55276 24464
rect 55316 24424 55317 24464
rect 55275 24415 55317 24424
rect 52971 23792 53013 23801
rect 52971 23752 52972 23792
rect 53012 23752 53013 23792
rect 52971 23743 53013 23752
rect 53643 23792 53685 23801
rect 53643 23752 53644 23792
rect 53684 23752 53685 23792
rect 53643 23743 53685 23752
rect 54795 23792 54837 23801
rect 54795 23752 54796 23792
rect 54836 23752 54837 23792
rect 54795 23743 54837 23752
rect 55084 23792 55124 23801
rect 55276 23792 55316 24415
rect 55372 24044 55412 24592
rect 55508 24592 55604 24632
rect 55468 24583 55508 24592
rect 55660 24548 55700 25927
rect 55755 25304 55797 25313
rect 55755 25264 55756 25304
rect 55796 25264 55797 25304
rect 55755 25255 55797 25264
rect 55948 25304 55988 26104
rect 56044 26095 56084 26104
rect 56332 26144 56372 26767
rect 56620 26732 56660 26741
rect 56428 26312 56468 26321
rect 56620 26312 56660 26692
rect 56468 26272 56660 26312
rect 56428 26263 56468 26272
rect 56332 26095 56372 26104
rect 56524 26144 56564 26153
rect 56524 25985 56564 26104
rect 56620 26144 56660 26153
rect 56523 25976 56565 25985
rect 56523 25936 56524 25976
rect 56564 25936 56565 25976
rect 56620 25976 56660 26104
rect 56812 26144 56852 27523
rect 56812 26095 56852 26104
rect 57004 26144 57044 26153
rect 56812 25976 56852 25985
rect 56620 25936 56812 25976
rect 56523 25927 56565 25936
rect 56812 25927 56852 25936
rect 57004 25313 57044 26104
rect 57100 26144 57140 26153
rect 55756 25170 55796 25255
rect 55852 25220 55892 25229
rect 55372 23995 55412 24004
rect 55564 24508 55700 24548
rect 55372 23792 55412 23801
rect 55276 23752 55372 23792
rect 52492 23668 52916 23708
rect 52299 23036 52341 23045
rect 52299 22996 52300 23036
rect 52340 22996 52341 23036
rect 52299 22987 52341 22996
rect 52011 22868 52053 22877
rect 52011 22828 52012 22868
rect 52052 22828 52053 22868
rect 52011 22819 52053 22828
rect 52012 22532 52052 22819
rect 52012 22483 52052 22492
rect 52107 22280 52149 22289
rect 52107 22240 52108 22280
rect 52148 22240 52149 22280
rect 52107 22231 52149 22240
rect 52300 22280 52340 22987
rect 52395 22784 52437 22793
rect 52395 22744 52396 22784
rect 52436 22744 52437 22784
rect 52395 22735 52437 22744
rect 52396 22532 52436 22735
rect 52396 22483 52436 22492
rect 52492 22280 52532 23668
rect 52972 23624 53012 23743
rect 54123 23708 54165 23717
rect 54123 23668 54124 23708
rect 54164 23668 54165 23708
rect 54123 23659 54165 23668
rect 52876 23584 53012 23624
rect 54124 23624 54164 23659
rect 54796 23658 54836 23743
rect 52876 23465 52916 23584
rect 54124 23573 54164 23584
rect 54892 23624 54932 23633
rect 52875 23456 52917 23465
rect 52875 23416 52876 23456
rect 52916 23416 52917 23456
rect 52875 23407 52917 23416
rect 52971 23372 53013 23381
rect 52971 23332 52972 23372
rect 53012 23332 53013 23372
rect 52971 23323 53013 23332
rect 52587 23288 52629 23297
rect 52587 23248 52588 23288
rect 52628 23248 52629 23288
rect 52587 23239 52629 23248
rect 52588 23120 52628 23239
rect 52684 23129 52724 23214
rect 52875 23204 52917 23213
rect 52875 23164 52876 23204
rect 52916 23164 52917 23204
rect 52875 23155 52917 23164
rect 52588 23071 52628 23080
rect 52683 23120 52725 23129
rect 52683 23080 52684 23120
rect 52724 23080 52725 23120
rect 52683 23071 52725 23080
rect 52779 22952 52821 22961
rect 52779 22912 52780 22952
rect 52820 22912 52821 22952
rect 52779 22903 52821 22912
rect 52684 22532 52724 22541
rect 52780 22532 52820 22903
rect 52724 22492 52820 22532
rect 52684 22289 52724 22492
rect 52588 22280 52628 22289
rect 52492 22240 52588 22280
rect 52108 22146 52148 22231
rect 52300 22205 52340 22240
rect 52299 22196 52341 22205
rect 52299 22156 52300 22196
rect 52340 22156 52341 22196
rect 52299 22147 52341 22156
rect 52588 21776 52628 22240
rect 52683 22280 52725 22289
rect 52683 22240 52684 22280
rect 52724 22240 52725 22280
rect 52683 22231 52725 22240
rect 52204 21736 52628 21776
rect 52012 19088 52052 19097
rect 52012 18509 52052 19048
rect 52011 18500 52053 18509
rect 52011 18460 52012 18500
rect 52052 18460 52053 18500
rect 52011 18451 52053 18460
rect 51916 18292 52148 18332
rect 51723 18283 51765 18292
rect 51628 16952 51668 16961
rect 51628 16232 51668 16241
rect 51532 16192 51628 16232
rect 51052 16064 51092 16073
rect 51052 15569 51092 16024
rect 51436 15905 51476 16192
rect 51435 15896 51477 15905
rect 51435 15856 51436 15896
rect 51476 15856 51477 15896
rect 51435 15847 51477 15856
rect 51628 15821 51668 16192
rect 51627 15812 51669 15821
rect 51627 15772 51628 15812
rect 51668 15772 51669 15812
rect 51627 15763 51669 15772
rect 51147 15644 51189 15653
rect 51147 15604 51148 15644
rect 51188 15604 51189 15644
rect 51147 15595 51189 15604
rect 50956 15392 50996 15520
rect 51051 15560 51093 15569
rect 51051 15520 51052 15560
rect 51092 15520 51093 15560
rect 51051 15511 51093 15520
rect 51148 15560 51188 15595
rect 51148 15509 51188 15520
rect 51532 15560 51572 15569
rect 50860 15352 50996 15392
rect 50764 14636 50804 14645
rect 50571 14384 50613 14393
rect 50571 14344 50572 14384
rect 50612 14344 50613 14384
rect 50571 14335 50613 14344
rect 50764 14225 50804 14596
rect 50763 14216 50805 14225
rect 50763 14176 50764 14216
rect 50804 14176 50805 14216
rect 50763 14167 50805 14176
rect 50860 13469 50900 15352
rect 51148 15308 51188 15317
rect 50956 15268 51148 15308
rect 50956 14888 50996 15268
rect 51148 15259 51188 15268
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 50956 14848 51284 14888
rect 51148 14720 51188 14729
rect 51052 14680 51148 14720
rect 50956 13880 50996 13889
rect 51052 13880 51092 14680
rect 51148 14671 51188 14680
rect 51244 14552 51284 14848
rect 51148 14512 51284 14552
rect 51148 14048 51188 14512
rect 51339 14216 51381 14225
rect 51339 14176 51340 14216
rect 51380 14176 51381 14216
rect 51339 14167 51381 14176
rect 51243 14132 51285 14141
rect 51243 14092 51244 14132
rect 51284 14092 51285 14132
rect 51243 14083 51285 14092
rect 51148 13999 51188 14008
rect 51244 14048 51284 14083
rect 51340 14082 51380 14167
rect 51244 13997 51284 14008
rect 51436 14048 51476 14057
rect 51532 14048 51572 15520
rect 51628 15560 51668 15569
rect 51628 14393 51668 15520
rect 51724 15560 51764 18283
rect 51915 17744 51957 17753
rect 51915 17704 51916 17744
rect 51956 17704 51957 17744
rect 51915 17695 51957 17704
rect 51820 16820 51860 16829
rect 51820 15905 51860 16780
rect 51819 15896 51861 15905
rect 51819 15856 51820 15896
rect 51860 15856 51861 15896
rect 51819 15847 51861 15856
rect 51627 14384 51669 14393
rect 51627 14344 51628 14384
rect 51668 14344 51669 14384
rect 51627 14335 51669 14344
rect 51476 14008 51572 14048
rect 51436 13999 51476 14008
rect 50996 13840 51092 13880
rect 50956 13831 50996 13840
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 50859 13460 50901 13469
rect 50859 13420 50860 13460
rect 50900 13420 50901 13460
rect 50859 13411 50901 13420
rect 51531 13460 51573 13469
rect 51531 13420 51532 13460
rect 51572 13420 51573 13460
rect 51531 13411 51573 13420
rect 50667 13208 50709 13217
rect 50667 13168 50668 13208
rect 50708 13168 50709 13208
rect 50667 13159 50709 13168
rect 50668 13074 50708 13159
rect 51532 12980 51572 13411
rect 51628 13301 51668 14335
rect 51627 13292 51669 13301
rect 51627 13252 51628 13292
rect 51668 13252 51669 13292
rect 51627 13243 51669 13252
rect 51724 13133 51764 15520
rect 51819 15560 51861 15569
rect 51819 15520 51820 15560
rect 51860 15520 51861 15560
rect 51819 15511 51861 15520
rect 51820 15426 51860 15511
rect 51819 13376 51861 13385
rect 51819 13336 51820 13376
rect 51860 13336 51861 13376
rect 51819 13327 51861 13336
rect 51723 13124 51765 13133
rect 51723 13084 51724 13124
rect 51764 13084 51765 13124
rect 51723 13075 51765 13084
rect 51532 12940 51668 12980
rect 50379 12872 50421 12881
rect 50379 12832 50380 12872
rect 50420 12832 50421 12872
rect 50379 12823 50421 12832
rect 50283 11948 50325 11957
rect 50283 11908 50284 11948
rect 50324 11908 50325 11948
rect 50283 11899 50325 11908
rect 50380 11789 50420 12823
rect 50955 12536 50997 12545
rect 50955 12496 50956 12536
rect 50996 12496 50997 12536
rect 50955 12487 50997 12496
rect 51628 12536 51668 12940
rect 51820 12713 51860 13327
rect 51916 12980 51956 17695
rect 52011 17324 52053 17333
rect 52011 17284 52012 17324
rect 52052 17284 52053 17324
rect 52011 17275 52053 17284
rect 52012 15989 52052 17275
rect 52011 15980 52053 15989
rect 52011 15940 52012 15980
rect 52052 15940 52053 15980
rect 52011 15931 52053 15940
rect 52011 15812 52053 15821
rect 52011 15772 52012 15812
rect 52052 15772 52053 15812
rect 52011 15763 52053 15772
rect 52012 14720 52052 15763
rect 52108 15392 52148 18292
rect 52204 17081 52244 21736
rect 52587 21608 52629 21617
rect 52587 21568 52588 21608
rect 52628 21568 52629 21608
rect 52587 21559 52629 21568
rect 52684 21608 52724 21617
rect 52876 21608 52916 23155
rect 52972 22037 53012 23323
rect 54315 23204 54357 23213
rect 54315 23164 54316 23204
rect 54356 23164 54357 23204
rect 54315 23155 54357 23164
rect 54316 23060 54356 23155
rect 54892 23060 54932 23584
rect 55084 23213 55124 23752
rect 55372 23743 55412 23752
rect 55564 23792 55604 24508
rect 55852 24464 55892 25180
rect 55948 24557 55988 25264
rect 57003 25304 57045 25313
rect 57003 25264 57004 25304
rect 57044 25264 57045 25304
rect 57003 25255 57045 25264
rect 57100 24725 57140 26104
rect 57099 24716 57141 24725
rect 57099 24676 57100 24716
rect 57140 24676 57141 24716
rect 57099 24667 57141 24676
rect 56331 24632 56373 24641
rect 56331 24592 56332 24632
rect 56372 24592 56373 24632
rect 56331 24583 56373 24592
rect 55947 24548 55989 24557
rect 55947 24508 55948 24548
rect 55988 24508 55989 24548
rect 55947 24499 55989 24508
rect 56332 24498 56372 24583
rect 55564 23743 55604 23752
rect 55660 24424 55892 24464
rect 55660 23792 55700 24424
rect 57196 23969 57236 29371
rect 57387 29168 57429 29177
rect 57387 29128 57388 29168
rect 57428 29128 57429 29168
rect 57387 29119 57429 29128
rect 57388 29034 57428 29119
rect 57291 27740 57333 27749
rect 57291 27700 57292 27740
rect 57332 27700 57333 27740
rect 57291 27691 57333 27700
rect 57292 27606 57332 27691
rect 57483 25976 57525 25985
rect 57483 25936 57484 25976
rect 57524 25936 57525 25976
rect 57483 25927 57525 25936
rect 57484 25304 57524 25927
rect 57484 25255 57524 25264
rect 57483 24548 57525 24557
rect 57483 24508 57484 24548
rect 57524 24508 57525 24548
rect 57483 24499 57525 24508
rect 57484 24414 57524 24499
rect 57195 23960 57237 23969
rect 57195 23920 57196 23960
rect 57236 23920 57237 23960
rect 57195 23911 57237 23920
rect 57580 23885 57620 29455
rect 58540 28916 58580 28925
rect 58540 28673 58580 28876
rect 58539 28664 58581 28673
rect 58539 28624 58540 28664
rect 58580 28624 58581 28664
rect 58539 28615 58581 28624
rect 59020 28580 59060 29871
rect 58828 28540 59060 28580
rect 57772 28496 57812 28505
rect 57676 28456 57772 28496
rect 57676 27656 57716 28456
rect 57772 28447 57812 28456
rect 57963 28160 58005 28169
rect 57963 28120 57964 28160
rect 58004 28120 58005 28160
rect 57963 28111 58005 28120
rect 58731 28160 58773 28169
rect 58731 28120 58732 28160
rect 58772 28120 58773 28160
rect 58731 28111 58773 28120
rect 57676 27607 57716 27616
rect 57964 26900 58004 28111
rect 58732 28026 58772 28111
rect 58540 27656 58580 27665
rect 58580 27616 58772 27656
rect 58540 27607 58580 27616
rect 58059 27320 58101 27329
rect 58059 27280 58060 27320
rect 58100 27280 58101 27320
rect 58059 27271 58101 27280
rect 57964 26851 58004 26860
rect 57675 26816 57717 26825
rect 57675 26776 57676 26816
rect 57716 26776 57717 26816
rect 57675 26767 57717 26776
rect 57676 26237 57716 26767
rect 58060 26741 58100 27271
rect 58539 27068 58581 27077
rect 58539 27028 58540 27068
rect 58580 27028 58581 27068
rect 58539 27019 58581 27028
rect 58155 26984 58197 26993
rect 58155 26944 58156 26984
rect 58196 26944 58197 26984
rect 58155 26935 58197 26944
rect 58156 26850 58196 26935
rect 58540 26934 58580 27019
rect 58347 26900 58389 26909
rect 58347 26860 58348 26900
rect 58388 26860 58389 26900
rect 58347 26851 58389 26860
rect 58348 26766 58388 26851
rect 58059 26732 58101 26741
rect 58059 26692 58060 26732
rect 58100 26692 58101 26732
rect 58059 26683 58101 26692
rect 57675 26228 57717 26237
rect 57675 26188 57676 26228
rect 57716 26188 57717 26228
rect 57675 26179 57717 26188
rect 57964 25976 58004 25985
rect 57868 25936 57964 25976
rect 57868 25304 57908 25936
rect 57964 25927 58004 25936
rect 57963 25808 58005 25817
rect 57963 25768 57964 25808
rect 58004 25768 58005 25808
rect 57963 25759 58005 25768
rect 57868 25255 57908 25264
rect 57675 24128 57717 24137
rect 57675 24088 57676 24128
rect 57716 24088 57717 24128
rect 57675 24079 57717 24088
rect 57579 23876 57621 23885
rect 57579 23836 57580 23876
rect 57620 23836 57621 23876
rect 57579 23827 57621 23836
rect 55660 23743 55700 23752
rect 55851 23792 55893 23801
rect 55851 23752 55852 23792
rect 55892 23752 55893 23792
rect 55851 23743 55893 23752
rect 56043 23792 56085 23801
rect 56043 23752 56044 23792
rect 56084 23752 56085 23792
rect 56043 23743 56085 23752
rect 56140 23792 56180 23801
rect 55852 23658 55892 23743
rect 55180 23624 55220 23633
rect 55948 23624 55988 23633
rect 55220 23584 55412 23624
rect 55180 23575 55220 23584
rect 55275 23456 55317 23465
rect 55275 23416 55276 23456
rect 55316 23416 55317 23456
rect 55275 23407 55317 23416
rect 55083 23204 55125 23213
rect 55083 23164 55084 23204
rect 55124 23164 55125 23204
rect 55083 23155 55125 23164
rect 54054 23036 54096 23045
rect 54054 22996 54055 23036
rect 54095 22996 54096 23036
rect 54316 23020 54385 23060
rect 54054 22987 54096 22996
rect 53544 22952 53586 22961
rect 53544 22912 53545 22952
rect 53585 22912 53586 22952
rect 53544 22903 53586 22912
rect 53545 22596 53585 22903
rect 53654 22868 53696 22877
rect 53654 22828 53655 22868
rect 53695 22828 53696 22868
rect 53654 22819 53696 22828
rect 53655 22596 53695 22819
rect 53944 22784 53986 22793
rect 53944 22744 53945 22784
rect 53985 22744 53986 22784
rect 53944 22735 53986 22744
rect 53945 22596 53985 22735
rect 54055 22596 54095 22987
rect 54345 22596 54385 23020
rect 54744 23036 54786 23045
rect 54744 22996 54745 23036
rect 54785 22996 54786 23036
rect 54892 23020 55185 23060
rect 54744 22987 54786 22996
rect 54454 22784 54496 22793
rect 54454 22744 54455 22784
rect 54495 22744 54496 22784
rect 54454 22735 54496 22744
rect 54455 22596 54495 22735
rect 54745 22596 54785 22987
rect 54854 22868 54896 22877
rect 54854 22828 54855 22868
rect 54895 22828 54896 22868
rect 54854 22819 54896 22828
rect 54855 22596 54895 22819
rect 55145 22596 55185 23020
rect 55276 22784 55316 23407
rect 55372 23060 55412 23584
rect 55659 23204 55701 23213
rect 55659 23164 55660 23204
rect 55700 23164 55701 23204
rect 55659 23155 55701 23164
rect 55660 23060 55700 23155
rect 55948 23060 55988 23584
rect 55372 23020 55585 23060
rect 55255 22744 55316 22784
rect 55255 22596 55295 22744
rect 55545 22596 55585 23020
rect 55655 23020 55700 23060
rect 55945 23020 55988 23060
rect 55655 22596 55695 23020
rect 55945 22596 55985 23020
rect 56044 22784 56084 23743
rect 56140 23549 56180 23752
rect 56428 23792 56468 23801
rect 56236 23624 56276 23633
rect 56139 23540 56181 23549
rect 56139 23500 56140 23540
rect 56180 23500 56181 23540
rect 56139 23491 56181 23500
rect 56236 23060 56276 23584
rect 56428 23297 56468 23752
rect 56811 23792 56853 23801
rect 56811 23752 56812 23792
rect 56852 23752 56853 23792
rect 56811 23743 56853 23752
rect 57291 23792 57333 23801
rect 57291 23752 57292 23792
rect 57332 23752 57333 23792
rect 57291 23743 57333 23752
rect 57676 23792 57716 24079
rect 57964 23792 58004 25759
rect 58060 25145 58100 26683
rect 58539 26648 58581 26657
rect 58539 26608 58540 26648
rect 58580 26608 58581 26648
rect 58539 26599 58581 26608
rect 58540 26514 58580 26599
rect 58348 26144 58388 26153
rect 58252 26104 58348 26144
rect 58155 25724 58197 25733
rect 58155 25684 58156 25724
rect 58196 25684 58197 25724
rect 58155 25675 58197 25684
rect 58059 25136 58101 25145
rect 58059 25096 58060 25136
rect 58100 25096 58101 25136
rect 58059 25087 58101 25096
rect 58059 24716 58101 24725
rect 58059 24676 58060 24716
rect 58100 24676 58101 24716
rect 58059 24667 58101 24676
rect 58060 24632 58100 24667
rect 58060 24581 58100 24592
rect 58156 24632 58196 25675
rect 58252 24800 58292 26104
rect 58348 26095 58388 26104
rect 58540 26144 58580 26153
rect 58540 25985 58580 26104
rect 58635 26144 58677 26153
rect 58635 26104 58636 26144
rect 58676 26104 58677 26144
rect 58635 26095 58677 26104
rect 58636 26010 58676 26095
rect 58347 25976 58389 25985
rect 58347 25936 58348 25976
rect 58388 25936 58389 25976
rect 58347 25927 58389 25936
rect 58539 25976 58581 25985
rect 58539 25936 58540 25976
rect 58580 25936 58581 25976
rect 58539 25927 58581 25936
rect 58348 25842 58388 25927
rect 58443 25892 58485 25901
rect 58443 25852 58444 25892
rect 58484 25852 58485 25892
rect 58443 25843 58485 25852
rect 58348 24800 58388 24809
rect 58252 24760 58348 24800
rect 58348 24751 58388 24760
rect 58156 24583 58196 24592
rect 58252 24632 58292 24641
rect 58444 24632 58484 25843
rect 58732 25304 58772 27616
rect 58828 27329 58868 28540
rect 59116 28496 59156 31723
rect 59692 31613 59732 32152
rect 59788 32152 59884 32192
rect 59691 31604 59733 31613
rect 59691 31564 59692 31604
rect 59732 31564 59733 31604
rect 59691 31555 59733 31564
rect 59788 31529 59828 32152
rect 59884 32143 59924 32152
rect 59980 32864 60020 34327
rect 60172 33797 60212 34411
rect 60364 34208 60404 34217
rect 60171 33788 60213 33797
rect 60171 33748 60172 33788
rect 60212 33748 60213 33788
rect 60171 33739 60213 33748
rect 60172 33140 60212 33739
rect 60364 33293 60404 34168
rect 60363 33284 60405 33293
rect 60363 33244 60364 33284
rect 60404 33244 60405 33284
rect 60363 33235 60405 33244
rect 60172 33100 60308 33140
rect 59884 31940 59924 31949
rect 59787 31520 59829 31529
rect 59787 31480 59788 31520
rect 59828 31480 59829 31520
rect 59787 31471 59829 31480
rect 59596 31352 59636 31361
rect 59212 31312 59596 31352
rect 59212 29840 59252 31312
rect 59596 31303 59636 31312
rect 59788 31352 59828 31361
rect 59692 31184 59732 31193
rect 59692 30773 59732 31144
rect 59691 30764 59733 30773
rect 59691 30724 59692 30764
rect 59732 30724 59733 30764
rect 59691 30715 59733 30724
rect 59691 30596 59733 30605
rect 59691 30556 59692 30596
rect 59732 30556 59733 30596
rect 59691 30547 59733 30556
rect 59307 30092 59349 30101
rect 59307 30052 59308 30092
rect 59348 30052 59349 30092
rect 59307 30043 59349 30052
rect 59212 29791 59252 29800
rect 59308 29840 59348 30043
rect 59403 30008 59445 30017
rect 59403 29968 59404 30008
rect 59444 29968 59445 30008
rect 59403 29959 59445 29968
rect 59308 29791 59348 29800
rect 59404 29840 59444 29959
rect 59404 29791 59444 29800
rect 59500 29840 59540 29851
rect 59500 29765 59540 29800
rect 59499 29756 59541 29765
rect 59499 29716 59500 29756
rect 59540 29716 59636 29756
rect 59499 29707 59541 29716
rect 59211 29588 59253 29597
rect 59211 29548 59212 29588
rect 59252 29548 59253 29588
rect 59211 29539 59253 29548
rect 59212 29084 59252 29539
rect 59596 29168 59636 29716
rect 59596 29119 59636 29128
rect 59692 29168 59732 30547
rect 59788 30269 59828 31312
rect 59884 31352 59924 31900
rect 59980 31697 60020 32824
rect 59979 31688 60021 31697
rect 59979 31648 59980 31688
rect 60020 31648 60021 31688
rect 59979 31639 60021 31648
rect 60075 31604 60117 31613
rect 60075 31564 60076 31604
rect 60116 31564 60117 31604
rect 60075 31555 60117 31564
rect 59979 31520 60021 31529
rect 59979 31480 59980 31520
rect 60020 31480 60021 31520
rect 59979 31471 60021 31480
rect 59884 31303 59924 31312
rect 59980 31184 60020 31471
rect 59884 31144 60020 31184
rect 59787 30260 59829 30269
rect 59787 30220 59788 30260
rect 59828 30220 59829 30260
rect 59787 30211 59829 30220
rect 59787 29840 59829 29849
rect 59787 29800 59788 29840
rect 59828 29800 59829 29840
rect 59787 29791 59829 29800
rect 59788 29706 59828 29791
rect 59884 29168 59924 31144
rect 60076 30689 60116 31555
rect 60075 30680 60117 30689
rect 60075 30640 60076 30680
rect 60116 30640 60117 30680
rect 60075 30631 60117 30640
rect 60172 30428 60212 30437
rect 60076 29840 60116 29849
rect 60076 29681 60116 29800
rect 60172 29840 60212 30388
rect 60172 29765 60212 29800
rect 60268 30428 60308 33100
rect 60364 32192 60404 32201
rect 60364 31277 60404 32152
rect 60460 31781 60500 36436
rect 60939 35888 60981 35897
rect 60939 35848 60940 35888
rect 60980 35848 60981 35888
rect 60939 35839 60981 35848
rect 60747 33032 60789 33041
rect 60747 32992 60748 33032
rect 60788 32992 60789 33032
rect 60747 32983 60789 32992
rect 60748 32192 60788 32983
rect 60748 32143 60788 32152
rect 60459 31772 60501 31781
rect 60459 31732 60460 31772
rect 60500 31732 60501 31772
rect 60459 31723 60501 31732
rect 60652 31436 60692 31445
rect 60459 31352 60501 31361
rect 60459 31312 60460 31352
rect 60500 31312 60501 31352
rect 60459 31303 60501 31312
rect 60363 31268 60405 31277
rect 60363 31228 60364 31268
rect 60404 31228 60405 31268
rect 60363 31219 60405 31228
rect 60460 31184 60500 31303
rect 60364 30428 60404 30437
rect 60268 30388 60364 30428
rect 60171 29756 60213 29765
rect 60171 29716 60172 29756
rect 60212 29716 60213 29756
rect 60171 29707 60213 29716
rect 60075 29672 60117 29681
rect 60172 29676 60212 29707
rect 60075 29632 60076 29672
rect 60116 29632 60117 29672
rect 60075 29623 60117 29632
rect 60268 29597 60308 30388
rect 60364 30379 60404 30388
rect 60460 30260 60500 31144
rect 60364 30220 60500 30260
rect 60556 30596 60596 30605
rect 60267 29588 60309 29597
rect 60267 29548 60268 29588
rect 60308 29548 60309 29588
rect 60267 29539 60309 29548
rect 59212 29035 59252 29044
rect 59404 29000 59444 29009
rect 59692 29000 59732 29128
rect 59444 28960 59732 29000
rect 59788 29128 59884 29168
rect 59404 28951 59444 28960
rect 59788 28748 59828 29128
rect 59884 29119 59924 29128
rect 60364 29168 60404 30220
rect 60556 30185 60596 30556
rect 60555 30176 60597 30185
rect 60555 30136 60556 30176
rect 60596 30136 60597 30176
rect 60555 30127 60597 30136
rect 60460 30008 60500 30017
rect 60460 29513 60500 29968
rect 60652 29924 60692 31396
rect 60940 30848 60980 35839
rect 61036 35216 61076 35225
rect 61036 34385 61076 35176
rect 61035 34376 61077 34385
rect 61035 34336 61036 34376
rect 61076 34336 61077 34376
rect 61035 34327 61077 34336
rect 61132 33545 61172 37939
rect 61900 37400 61940 38032
rect 63531 37988 63573 37997
rect 63531 37948 63532 37988
rect 63572 37948 63573 37988
rect 63531 37939 63573 37948
rect 63532 37854 63572 37939
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 62092 37400 62132 37409
rect 61900 37360 62092 37400
rect 62092 37351 62132 37360
rect 62955 37400 62997 37409
rect 62955 37360 62956 37400
rect 62996 37360 62997 37400
rect 62955 37351 62997 37360
rect 61611 37316 61653 37325
rect 61611 37276 61612 37316
rect 61652 37276 61653 37316
rect 61611 37267 61653 37276
rect 61708 37316 61748 37325
rect 61748 37276 62036 37316
rect 61708 37267 61748 37276
rect 61516 37232 61556 37241
rect 61516 36989 61556 37192
rect 61515 36980 61557 36989
rect 61515 36940 61516 36980
rect 61556 36940 61557 36980
rect 61515 36931 61557 36940
rect 61419 36728 61461 36737
rect 61419 36688 61420 36728
rect 61460 36688 61461 36728
rect 61419 36679 61461 36688
rect 61516 36728 61556 36737
rect 61420 36594 61460 36679
rect 61516 36224 61556 36688
rect 61228 36184 61556 36224
rect 61612 36728 61652 37267
rect 61996 36896 62036 37276
rect 62956 37266 62996 37351
rect 63435 37316 63477 37325
rect 63435 37276 63436 37316
rect 63476 37276 63477 37316
rect 63435 37267 63477 37276
rect 61996 36847 62036 36856
rect 61228 35897 61268 36184
rect 61419 36056 61461 36065
rect 61419 36016 61420 36056
rect 61460 36016 61461 36056
rect 61612 36056 61652 36688
rect 61708 36728 61748 36737
rect 61900 36728 61940 36737
rect 61748 36688 61900 36728
rect 61708 36679 61748 36688
rect 61900 36679 61940 36688
rect 62092 36728 62132 36737
rect 62092 36569 62132 36688
rect 62188 36728 62228 36737
rect 63148 36728 63188 36737
rect 62091 36560 62133 36569
rect 62091 36520 62092 36560
rect 62132 36520 62133 36560
rect 62091 36511 62133 36520
rect 62188 36065 62228 36688
rect 62956 36688 63148 36728
rect 62187 36056 62229 36065
rect 61612 36016 61940 36056
rect 61419 36007 61461 36016
rect 61227 35888 61269 35897
rect 61227 35848 61228 35888
rect 61268 35848 61269 35888
rect 61227 35839 61269 35848
rect 61324 35888 61364 35897
rect 61324 33629 61364 35848
rect 61420 35804 61460 36007
rect 61516 35981 61556 36012
rect 61515 35972 61557 35981
rect 61515 35932 61516 35972
rect 61556 35932 61557 35972
rect 61515 35923 61557 35932
rect 61420 35755 61460 35764
rect 61516 35888 61556 35923
rect 61419 35552 61461 35561
rect 61419 35512 61420 35552
rect 61460 35512 61461 35552
rect 61419 35503 61461 35512
rect 61420 35057 61460 35503
rect 61419 35048 61461 35057
rect 61419 35008 61420 35048
rect 61460 35008 61461 35048
rect 61419 34999 61461 35008
rect 61323 33620 61365 33629
rect 61323 33580 61324 33620
rect 61364 33580 61365 33620
rect 61323 33571 61365 33580
rect 61131 33536 61173 33545
rect 61131 33496 61132 33536
rect 61172 33496 61173 33536
rect 61131 33487 61173 33496
rect 61323 33032 61365 33041
rect 61323 32992 61324 33032
rect 61364 32992 61365 33032
rect 61323 32983 61365 32992
rect 61324 32898 61364 32983
rect 61132 32696 61172 32705
rect 61132 31865 61172 32656
rect 61131 31856 61173 31865
rect 61131 31816 61132 31856
rect 61172 31816 61173 31856
rect 61131 31807 61173 31816
rect 61132 31520 61172 31529
rect 60940 30799 60980 30808
rect 61036 31480 61132 31520
rect 60747 30596 60789 30605
rect 60747 30556 60748 30596
rect 60788 30556 60789 30596
rect 60747 30547 60789 30556
rect 60748 30462 60788 30547
rect 60940 30437 60980 30522
rect 60939 30428 60981 30437
rect 60939 30388 60940 30428
rect 60980 30388 60981 30428
rect 60939 30379 60981 30388
rect 60939 30260 60981 30269
rect 60939 30220 60940 30260
rect 60980 30220 60981 30260
rect 60939 30211 60981 30220
rect 60652 29884 60788 29924
rect 60652 29756 60692 29765
rect 60459 29504 60501 29513
rect 60459 29464 60460 29504
rect 60500 29464 60501 29504
rect 60459 29455 60501 29464
rect 60460 29336 60500 29345
rect 60652 29336 60692 29716
rect 60500 29296 60692 29336
rect 60460 29287 60500 29296
rect 60364 29119 60404 29128
rect 60556 29168 60596 29179
rect 60556 29093 60596 29128
rect 60651 29168 60693 29177
rect 60651 29128 60652 29168
rect 60692 29128 60693 29168
rect 60651 29119 60693 29128
rect 60555 29084 60597 29093
rect 60555 29044 60556 29084
rect 60596 29044 60597 29084
rect 60555 29035 60597 29044
rect 60652 29034 60692 29119
rect 59884 28916 59924 28925
rect 59924 28876 60116 28916
rect 59884 28867 59924 28876
rect 59788 28708 59924 28748
rect 59020 28456 59156 28496
rect 59307 28496 59349 28505
rect 59307 28456 59308 28496
rect 59348 28456 59349 28496
rect 58924 28412 58964 28421
rect 58924 28085 58964 28372
rect 58923 28076 58965 28085
rect 58923 28036 58924 28076
rect 58964 28036 58965 28076
rect 58923 28027 58965 28036
rect 58827 27320 58869 27329
rect 58827 27280 58828 27320
rect 58868 27280 58869 27320
rect 58827 27271 58869 27280
rect 59020 27161 59060 28456
rect 59307 28447 59349 28456
rect 59115 28328 59157 28337
rect 59115 28288 59116 28328
rect 59156 28288 59157 28328
rect 59115 28279 59157 28288
rect 59212 28328 59252 28337
rect 59019 27152 59061 27161
rect 59019 27112 59020 27152
rect 59060 27112 59061 27152
rect 59019 27103 59061 27112
rect 58827 26984 58869 26993
rect 58827 26944 58828 26984
rect 58868 26944 58869 26984
rect 58827 26935 58869 26944
rect 58828 26816 58868 26935
rect 58828 26767 58868 26776
rect 59019 26816 59061 26825
rect 59019 26776 59020 26816
rect 59060 26776 59061 26816
rect 59019 26767 59061 26776
rect 59116 26816 59156 28279
rect 59212 26993 59252 28288
rect 59308 28328 59348 28447
rect 59211 26984 59253 26993
rect 59211 26944 59212 26984
rect 59252 26944 59253 26984
rect 59211 26935 59253 26944
rect 59116 26767 59156 26776
rect 59020 26682 59060 26767
rect 58827 26648 58869 26657
rect 58827 26608 58828 26648
rect 58868 26608 58869 26648
rect 58827 26599 58869 26608
rect 58924 26648 58964 26657
rect 58828 26060 58868 26599
rect 58924 26153 58964 26608
rect 59020 26312 59060 26321
rect 59212 26312 59252 26935
rect 59308 26564 59348 28288
rect 59596 28412 59636 28421
rect 59404 28160 59444 28169
rect 59404 27656 59444 28120
rect 59596 27833 59636 28372
rect 59691 28328 59733 28337
rect 59691 28288 59692 28328
rect 59732 28288 59733 28328
rect 59691 28279 59733 28288
rect 59595 27824 59637 27833
rect 59595 27784 59596 27824
rect 59636 27784 59637 27824
rect 59595 27775 59637 27784
rect 59692 27824 59732 28279
rect 59788 28160 59828 28171
rect 59884 28169 59924 28708
rect 59788 28085 59828 28120
rect 59883 28160 59925 28169
rect 59883 28120 59884 28160
rect 59924 28120 59925 28160
rect 60076 28160 60116 28876
rect 60748 28832 60788 29884
rect 60843 29504 60885 29513
rect 60843 29464 60844 29504
rect 60884 29464 60885 29504
rect 60843 29455 60885 29464
rect 60844 29168 60884 29455
rect 60844 29119 60884 29128
rect 60940 29252 60980 30211
rect 61036 29840 61076 31480
rect 61132 31471 61172 31480
rect 61131 30680 61173 30689
rect 61131 30640 61132 30680
rect 61172 30640 61173 30680
rect 61131 30631 61173 30640
rect 61324 30680 61364 30689
rect 61132 30546 61172 30631
rect 61228 30428 61268 30437
rect 61131 30176 61173 30185
rect 61131 30136 61132 30176
rect 61172 30136 61173 30176
rect 61131 30127 61173 30136
rect 61036 29791 61076 29800
rect 60940 29093 60980 29212
rect 61035 29252 61077 29261
rect 61035 29212 61036 29252
rect 61076 29212 61077 29252
rect 61035 29203 61077 29212
rect 61036 29168 61076 29203
rect 61036 29117 61076 29128
rect 60939 29084 60981 29093
rect 60939 29044 60940 29084
rect 60980 29044 60981 29084
rect 60939 29035 60981 29044
rect 60748 28792 60980 28832
rect 60843 28580 60885 28589
rect 60843 28540 60844 28580
rect 60884 28540 60885 28580
rect 60843 28531 60885 28540
rect 60172 28337 60212 28422
rect 60171 28328 60213 28337
rect 60171 28288 60172 28328
rect 60212 28288 60213 28328
rect 60171 28279 60213 28288
rect 60363 28328 60405 28337
rect 60363 28288 60364 28328
rect 60404 28288 60405 28328
rect 60363 28279 60405 28288
rect 60460 28328 60500 28337
rect 60268 28160 60308 28169
rect 60076 28120 60212 28160
rect 59883 28111 59925 28120
rect 59787 28076 59829 28085
rect 59787 28036 59788 28076
rect 59828 28036 59829 28076
rect 59787 28027 59829 28036
rect 59884 27833 59924 28111
rect 60075 27908 60117 27917
rect 60075 27868 60076 27908
rect 60116 27868 60117 27908
rect 60075 27859 60117 27868
rect 59692 27775 59732 27784
rect 59883 27824 59925 27833
rect 59883 27784 59884 27824
rect 59924 27784 59925 27824
rect 59883 27775 59925 27784
rect 59979 27740 60021 27749
rect 59979 27700 59980 27740
rect 60020 27700 60021 27740
rect 59979 27691 60021 27700
rect 59884 27656 59924 27665
rect 59404 27616 59884 27656
rect 59884 27607 59924 27616
rect 59980 27606 60020 27691
rect 60076 27656 60116 27859
rect 60076 27607 60116 27616
rect 60172 27656 60212 28120
rect 60268 27740 60308 28120
rect 60364 27917 60404 28279
rect 60460 28085 60500 28288
rect 60652 28328 60692 28337
rect 60459 28076 60501 28085
rect 60459 28036 60460 28076
rect 60500 28036 60501 28076
rect 60459 28027 60501 28036
rect 60363 27908 60405 27917
rect 60363 27868 60364 27908
rect 60404 27868 60405 27908
rect 60363 27859 60405 27868
rect 60556 27740 60596 27749
rect 60268 27700 60556 27740
rect 60556 27691 60596 27700
rect 60172 27607 60212 27616
rect 60652 27497 60692 28288
rect 60747 28328 60789 28337
rect 60747 28288 60748 28328
rect 60788 28288 60789 28328
rect 60747 28279 60789 28288
rect 60844 28328 60884 28531
rect 60940 28412 60980 28792
rect 61036 28580 61076 28589
rect 61132 28580 61172 30127
rect 61228 29177 61268 30388
rect 61324 29681 61364 30640
rect 61420 29933 61460 34999
rect 61516 34880 61556 35848
rect 61611 35888 61653 35897
rect 61611 35848 61612 35888
rect 61652 35848 61653 35888
rect 61611 35839 61653 35848
rect 61612 35754 61652 35839
rect 61708 35561 61748 36016
rect 61900 35888 61940 36016
rect 62187 36016 62188 36056
rect 62228 36016 62229 36056
rect 62187 36007 62229 36016
rect 61900 35839 61940 35848
rect 61996 35888 62036 35899
rect 61996 35813 62036 35848
rect 62091 35888 62133 35897
rect 62091 35848 62092 35888
rect 62132 35848 62133 35888
rect 62091 35839 62133 35848
rect 62667 35888 62709 35897
rect 62667 35848 62668 35888
rect 62708 35848 62709 35888
rect 62667 35839 62709 35848
rect 61995 35804 62037 35813
rect 61995 35764 61996 35804
rect 62036 35764 62037 35804
rect 61995 35755 62037 35764
rect 62092 35754 62132 35839
rect 61804 35720 61844 35729
rect 61707 35552 61749 35561
rect 61707 35512 61708 35552
rect 61748 35512 61749 35552
rect 61707 35503 61749 35512
rect 61516 34840 61652 34880
rect 61515 34712 61557 34721
rect 61515 34672 61516 34712
rect 61556 34672 61557 34712
rect 61515 34663 61557 34672
rect 61516 33140 61556 34663
rect 61612 33713 61652 34840
rect 61804 34376 61844 35680
rect 62668 35300 62708 35839
rect 62188 34964 62228 34973
rect 62188 34805 62228 34924
rect 62380 34964 62420 34973
rect 62187 34796 62229 34805
rect 62187 34756 62188 34796
rect 62228 34756 62229 34796
rect 62187 34747 62229 34756
rect 61900 34553 61940 34638
rect 61899 34544 61941 34553
rect 61899 34504 61900 34544
rect 61940 34504 61941 34544
rect 61899 34495 61941 34504
rect 61900 34376 61940 34385
rect 61804 34336 61900 34376
rect 61900 34327 61940 34336
rect 62091 34376 62133 34385
rect 62091 34336 62092 34376
rect 62132 34336 62133 34376
rect 62091 34327 62133 34336
rect 62188 34376 62228 34385
rect 62228 34336 62324 34376
rect 62188 34327 62228 34336
rect 62092 34242 62132 34327
rect 62091 34040 62133 34049
rect 62091 34000 62092 34040
rect 62132 34000 62133 34040
rect 62091 33991 62133 34000
rect 61611 33704 61653 33713
rect 61611 33664 61612 33704
rect 61652 33664 61653 33704
rect 61611 33655 61653 33664
rect 61516 33100 61844 33140
rect 61515 33032 61557 33041
rect 61515 32992 61516 33032
rect 61556 32992 61557 33032
rect 61515 32983 61557 32992
rect 61516 31856 61556 32983
rect 61612 32192 61652 32203
rect 61612 32117 61652 32152
rect 61611 32108 61653 32117
rect 61611 32068 61612 32108
rect 61652 32068 61653 32108
rect 61611 32059 61653 32068
rect 61516 31816 61748 31856
rect 61708 30848 61748 31816
rect 61708 30799 61748 30808
rect 61516 30596 61556 30605
rect 61804 30596 61844 33100
rect 61899 32108 61941 32117
rect 61899 32068 61900 32108
rect 61940 32068 61941 32108
rect 61899 32059 61941 32068
rect 61900 31697 61940 32059
rect 61899 31688 61941 31697
rect 61899 31648 61900 31688
rect 61940 31648 61941 31688
rect 61899 31639 61941 31648
rect 61556 30556 61844 30596
rect 61419 29924 61461 29933
rect 61419 29884 61420 29924
rect 61460 29884 61461 29924
rect 61419 29875 61461 29884
rect 61323 29672 61365 29681
rect 61323 29632 61324 29672
rect 61364 29632 61365 29672
rect 61323 29623 61365 29632
rect 61227 29168 61269 29177
rect 61227 29128 61228 29168
rect 61268 29128 61269 29168
rect 61227 29119 61269 29128
rect 61516 28589 61556 30556
rect 61708 30428 61748 30437
rect 61611 29504 61653 29513
rect 61611 29464 61612 29504
rect 61652 29464 61653 29504
rect 61611 29455 61653 29464
rect 61076 28540 61172 28580
rect 61515 28580 61557 28589
rect 61515 28540 61516 28580
rect 61556 28540 61557 28580
rect 61036 28531 61076 28540
rect 61515 28531 61557 28540
rect 61612 28580 61652 29455
rect 61708 29261 61748 30388
rect 61900 29840 61940 31639
rect 62092 31361 62132 33991
rect 62284 33788 62324 34336
rect 62380 33872 62420 34924
rect 62668 34805 62708 35260
rect 62764 35216 62804 35225
rect 62667 34796 62709 34805
rect 62667 34756 62668 34796
rect 62708 34756 62709 34796
rect 62667 34747 62709 34756
rect 62764 34628 62804 35176
rect 62668 34588 62804 34628
rect 62956 35216 62996 36688
rect 63148 36679 63188 36688
rect 63436 36728 63476 37267
rect 63531 37232 63573 37241
rect 63531 37192 63532 37232
rect 63572 37192 63573 37232
rect 63531 37183 63573 37192
rect 63532 36812 63572 37183
rect 63532 36737 63572 36772
rect 63436 36679 63476 36688
rect 63531 36728 63573 36737
rect 63531 36688 63532 36728
rect 63572 36688 63573 36728
rect 63531 36679 63573 36688
rect 63532 36648 63572 36679
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 63052 35216 63092 35225
rect 62956 35176 63052 35216
rect 62571 34544 62613 34553
rect 62571 34504 62572 34544
rect 62612 34504 62613 34544
rect 62571 34495 62613 34504
rect 62572 34376 62612 34495
rect 62668 34469 62708 34588
rect 62667 34460 62709 34469
rect 62667 34420 62668 34460
rect 62708 34420 62709 34460
rect 62667 34411 62709 34420
rect 62764 34385 62804 34470
rect 62572 34049 62612 34336
rect 62763 34376 62805 34385
rect 62763 34336 62764 34376
rect 62804 34336 62805 34376
rect 62763 34327 62805 34336
rect 62860 34376 62900 34385
rect 62667 34292 62709 34301
rect 62667 34252 62668 34292
rect 62708 34252 62709 34292
rect 62667 34243 62709 34252
rect 62668 34158 62708 34243
rect 62571 34040 62613 34049
rect 62571 34000 62572 34040
rect 62612 34000 62613 34040
rect 62571 33991 62613 34000
rect 62380 33832 62708 33872
rect 62284 33739 62324 33748
rect 62188 33704 62228 33715
rect 62188 33629 62228 33664
rect 62379 33704 62421 33713
rect 62379 33664 62380 33704
rect 62420 33664 62421 33704
rect 62379 33655 62421 33664
rect 62476 33704 62516 33713
rect 62668 33704 62708 33832
rect 62764 33788 62804 34327
rect 62860 34049 62900 34336
rect 62859 34040 62901 34049
rect 62859 34000 62860 34040
rect 62900 34000 62901 34040
rect 62859 33991 62901 34000
rect 62764 33739 62804 33748
rect 62516 33664 62612 33704
rect 62476 33655 62516 33664
rect 62187 33620 62229 33629
rect 62187 33580 62188 33620
rect 62228 33580 62229 33620
rect 62187 33571 62229 33580
rect 62091 31352 62133 31361
rect 62091 31312 62092 31352
rect 62132 31312 62133 31352
rect 62091 31303 62133 31312
rect 62188 30428 62228 33571
rect 62380 33570 62420 33655
rect 62475 33536 62517 33545
rect 62475 33496 62476 33536
rect 62516 33496 62517 33536
rect 62475 33487 62517 33496
rect 62476 32957 62516 33487
rect 62572 33116 62612 33664
rect 62668 33655 62708 33664
rect 62860 33704 62900 33713
rect 62860 33125 62900 33664
rect 62956 33140 62996 35176
rect 63052 35167 63092 35176
rect 63532 35048 63572 35057
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 63243 34460 63285 34469
rect 63243 34420 63244 34460
rect 63284 34420 63285 34460
rect 63243 34411 63285 34420
rect 63051 34292 63093 34301
rect 63051 34252 63052 34292
rect 63092 34252 63093 34292
rect 63051 34243 63093 34252
rect 63052 34158 63092 34243
rect 63244 34133 63284 34411
rect 63436 34376 63476 34385
rect 63532 34376 63572 35008
rect 63628 34469 63668 38200
rect 63724 36569 63764 38200
rect 63820 38240 63860 38368
rect 64108 38324 64148 38368
rect 64108 38275 64148 38284
rect 70155 38324 70197 38333
rect 70155 38284 70156 38324
rect 70196 38284 70197 38324
rect 70155 38275 70197 38284
rect 71403 38324 71445 38333
rect 71403 38284 71404 38324
rect 71444 38284 71445 38324
rect 71403 38275 71445 38284
rect 63820 38191 63860 38200
rect 64012 38240 64052 38249
rect 64012 37460 64052 38200
rect 63916 37420 64052 37460
rect 64204 38240 64244 38249
rect 63819 36728 63861 36737
rect 63819 36688 63820 36728
rect 63860 36688 63861 36728
rect 63819 36679 63861 36688
rect 63723 36560 63765 36569
rect 63723 36520 63724 36560
rect 63764 36520 63765 36560
rect 63723 36511 63765 36520
rect 63820 36560 63860 36679
rect 63916 36644 63956 37420
rect 64204 37325 64244 38200
rect 67467 38240 67509 38249
rect 68044 38240 68084 38249
rect 67467 38200 67468 38240
rect 67508 38200 67509 38240
rect 67467 38191 67509 38200
rect 67948 38200 68044 38240
rect 64588 38072 64628 38081
rect 64299 37988 64341 37997
rect 64299 37948 64300 37988
rect 64340 37948 64341 37988
rect 64299 37939 64341 37948
rect 64300 37400 64340 37939
rect 64588 37460 64628 38032
rect 66220 38072 66260 38081
rect 66220 37460 66260 38032
rect 64588 37420 64724 37460
rect 64300 37351 64340 37360
rect 64684 37400 64724 37420
rect 66124 37420 66260 37460
rect 64684 37351 64724 37360
rect 65547 37400 65589 37409
rect 65547 37360 65548 37400
rect 65588 37360 65589 37400
rect 65547 37351 65589 37360
rect 64203 37316 64245 37325
rect 64203 37276 64204 37316
rect 64244 37276 64245 37316
rect 64203 37267 64245 37276
rect 64107 37232 64149 37241
rect 64107 37192 64108 37232
rect 64148 37192 64149 37232
rect 64107 37183 64149 37192
rect 64108 37098 64148 37183
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 65548 36737 65588 37351
rect 64011 36728 64053 36737
rect 64011 36688 64012 36728
rect 64052 36688 64053 36728
rect 64011 36679 64053 36688
rect 64204 36728 64244 36737
rect 63915 36604 63956 36644
rect 63915 36560 63955 36604
rect 64012 36594 64052 36679
rect 64107 36560 64149 36569
rect 63915 36520 63956 36560
rect 63820 36511 63860 36520
rect 63627 34460 63669 34469
rect 63627 34420 63628 34460
rect 63668 34420 63669 34460
rect 63627 34411 63669 34420
rect 63476 34336 63572 34376
rect 63436 34327 63476 34336
rect 63243 34124 63285 34133
rect 63243 34084 63244 34124
rect 63284 34084 63285 34124
rect 63243 34075 63285 34084
rect 63147 34040 63189 34049
rect 63147 34000 63148 34040
rect 63188 34000 63189 34040
rect 63147 33991 63189 34000
rect 63051 33788 63093 33797
rect 63051 33748 63052 33788
rect 63092 33748 63093 33788
rect 63051 33739 63093 33748
rect 63148 33788 63188 33991
rect 63148 33739 63188 33748
rect 63052 33704 63092 33739
rect 63052 33653 63092 33664
rect 63244 33704 63284 34075
rect 63244 33655 63284 33664
rect 63724 33536 63764 33545
rect 63628 33496 63724 33536
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 62859 33116 62901 33125
rect 62572 33076 62708 33116
rect 62475 32948 62517 32957
rect 62475 32908 62476 32948
rect 62516 32908 62517 32948
rect 62475 32899 62517 32908
rect 62283 32864 62325 32873
rect 62283 32824 62284 32864
rect 62324 32824 62325 32864
rect 62283 32815 62325 32824
rect 62476 32864 62516 32899
rect 62572 32873 62612 32958
rect 62284 30605 62324 32815
rect 62476 32814 62516 32824
rect 62571 32864 62613 32873
rect 62571 32824 62572 32864
rect 62612 32824 62613 32864
rect 62571 32815 62613 32824
rect 62668 32864 62708 33076
rect 62859 33076 62860 33116
rect 62900 33076 62901 33116
rect 62956 33100 63092 33140
rect 62859 33067 62901 33076
rect 62380 32696 62420 32705
rect 62420 32656 62612 32696
rect 62380 32647 62420 32656
rect 62475 32108 62517 32117
rect 62475 32068 62476 32108
rect 62516 32068 62517 32108
rect 62475 32059 62517 32068
rect 62476 30689 62516 32059
rect 62572 31352 62612 32656
rect 62668 32537 62708 32824
rect 62667 32528 62709 32537
rect 62667 32488 62668 32528
rect 62708 32488 62709 32528
rect 62667 32479 62709 32488
rect 62668 32360 62708 32479
rect 62764 32360 62804 32369
rect 62668 32320 62764 32360
rect 62764 32311 62804 32320
rect 63052 32285 63092 33100
rect 63628 32864 63668 33496
rect 63724 33487 63764 33496
rect 63916 33140 63956 36520
rect 64107 36520 64108 36560
rect 64148 36520 64149 36560
rect 64107 36511 64149 36520
rect 64108 36426 64148 36511
rect 64204 35972 64244 36688
rect 65547 36728 65589 36737
rect 65547 36688 65548 36728
rect 65588 36688 65589 36728
rect 65547 36679 65589 36688
rect 65740 36728 65780 36737
rect 64108 35932 64244 35972
rect 64108 34721 64148 35932
rect 64588 35888 64628 35897
rect 65452 35888 65492 35897
rect 65548 35888 65588 36679
rect 65740 36485 65780 36688
rect 66124 36728 66164 37420
rect 66315 37400 66357 37409
rect 66315 37360 66316 37400
rect 66356 37360 66357 37400
rect 66315 37351 66357 37360
rect 67084 37400 67124 37409
rect 66124 36679 66164 36688
rect 65739 36476 65781 36485
rect 65739 36436 65740 36476
rect 65780 36436 65781 36476
rect 65739 36427 65781 36436
rect 64628 35848 64820 35888
rect 64588 35839 64628 35848
rect 64203 35804 64245 35813
rect 64203 35764 64204 35804
rect 64244 35764 64245 35804
rect 64203 35755 64245 35764
rect 64204 35670 64244 35755
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 64684 35048 64724 35057
rect 64780 35048 64820 35848
rect 65492 35848 65588 35888
rect 65452 35839 65492 35848
rect 66027 35720 66069 35729
rect 66027 35680 66028 35720
rect 66068 35680 66069 35720
rect 66027 35671 66069 35680
rect 65163 35636 65205 35645
rect 65163 35596 65164 35636
rect 65204 35596 65205 35636
rect 65163 35587 65205 35596
rect 64724 35008 64820 35048
rect 64684 34999 64724 35008
rect 64107 34712 64149 34721
rect 64107 34672 64108 34712
rect 64148 34672 64149 34712
rect 64107 34663 64149 34672
rect 64300 34376 64340 34385
rect 63628 32815 63668 32824
rect 63724 33100 63956 33140
rect 64204 34336 64300 34376
rect 64107 33116 64149 33125
rect 63244 32780 63284 32789
rect 63148 32740 63244 32780
rect 63051 32276 63093 32285
rect 63051 32236 63052 32276
rect 63092 32236 63093 32276
rect 63051 32227 63093 32236
rect 63052 32192 63092 32227
rect 63052 32142 63092 32152
rect 62859 31940 62901 31949
rect 63148 31940 63188 32740
rect 63244 32731 63284 32740
rect 63724 32696 63764 33100
rect 64107 33076 64108 33116
rect 64148 33076 64149 33116
rect 64107 33067 64149 33076
rect 64011 32948 64053 32957
rect 64011 32908 64012 32948
rect 64052 32908 64053 32948
rect 64011 32899 64053 32908
rect 63628 32656 63764 32696
rect 63435 32528 63477 32537
rect 63435 32488 63436 32528
rect 63476 32488 63477 32528
rect 63435 32479 63477 32488
rect 63243 32276 63285 32285
rect 63436 32276 63476 32479
rect 63243 32236 63244 32276
rect 63284 32236 63380 32276
rect 63243 32227 63285 32236
rect 63340 32219 63380 32236
rect 63436 32227 63476 32236
rect 63340 32170 63380 32179
rect 62859 31900 62860 31940
rect 62900 31900 62901 31940
rect 62859 31891 62901 31900
rect 62956 31900 63188 31940
rect 63531 31940 63573 31949
rect 63531 31900 63532 31940
rect 63572 31900 63573 31940
rect 62860 31772 62900 31891
rect 62572 31303 62612 31312
rect 62764 31732 62900 31772
rect 62764 31352 62804 31732
rect 62956 31604 62996 31900
rect 63531 31891 63573 31900
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 63052 31604 63092 31613
rect 63532 31604 63572 31891
rect 63628 31856 63668 32656
rect 63916 32192 63956 32201
rect 63724 32024 63764 32033
rect 63916 32024 63956 32152
rect 64012 32108 64052 32899
rect 64108 32285 64148 33067
rect 64204 32864 64244 34336
rect 64300 34327 64340 34336
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 65164 33140 65204 35587
rect 65835 35384 65877 35393
rect 65835 35344 65836 35384
rect 65876 35344 65877 35384
rect 65835 35335 65877 35344
rect 65836 35250 65876 35335
rect 65932 35216 65972 35225
rect 65932 35057 65972 35176
rect 66028 35216 66068 35671
rect 65931 35048 65973 35057
rect 65931 35008 65932 35048
rect 65972 35008 65973 35048
rect 65931 34999 65973 35008
rect 65452 34208 65492 34219
rect 65452 34133 65492 34168
rect 65451 34124 65493 34133
rect 65451 34084 65452 34124
rect 65492 34084 65493 34124
rect 65451 34075 65493 34084
rect 65932 33545 65972 34999
rect 65931 33536 65973 33545
rect 65931 33496 65932 33536
rect 65972 33496 65973 33536
rect 65931 33487 65973 33496
rect 66028 33452 66068 35176
rect 66123 35216 66165 35225
rect 66123 35176 66124 35216
rect 66164 35176 66165 35216
rect 66123 35167 66165 35176
rect 66124 35082 66164 35167
rect 66124 34376 66164 34385
rect 66124 33629 66164 34336
rect 66316 34376 66356 37351
rect 66700 37325 66740 37356
rect 66699 37316 66741 37325
rect 66699 37276 66700 37316
rect 66740 37276 66741 37316
rect 66699 37267 66741 37276
rect 66700 37232 66740 37267
rect 66700 35981 66740 37192
rect 66987 36728 67029 36737
rect 66987 36688 66988 36728
rect 67028 36688 67029 36728
rect 66987 36679 67029 36688
rect 66988 36594 67028 36679
rect 67084 36233 67124 37360
rect 67275 37400 67317 37409
rect 67275 37360 67276 37400
rect 67316 37360 67317 37400
rect 67275 37351 67317 37360
rect 67372 37400 67412 37409
rect 67276 37266 67316 37351
rect 67180 37232 67220 37241
rect 67083 36224 67125 36233
rect 67083 36184 67084 36224
rect 67124 36184 67125 36224
rect 67083 36175 67125 36184
rect 66699 35972 66741 35981
rect 66699 35932 66700 35972
rect 66740 35932 66741 35972
rect 66699 35923 66741 35932
rect 66796 35888 66836 35897
rect 66604 35720 66644 35729
rect 66604 35225 66644 35680
rect 66796 35393 66836 35848
rect 66987 35888 67029 35897
rect 66987 35848 66988 35888
rect 67028 35848 67029 35888
rect 66987 35839 67029 35848
rect 67084 35888 67124 35897
rect 67180 35888 67220 37192
rect 67372 36905 67412 37360
rect 67371 36896 67413 36905
rect 67371 36856 67372 36896
rect 67412 36856 67413 36896
rect 67371 36847 67413 36856
rect 67468 36056 67508 38191
rect 67852 38156 67892 38165
rect 67755 38072 67797 38081
rect 67852 38072 67892 38116
rect 67755 38032 67756 38072
rect 67796 38032 67892 38072
rect 67755 38023 67797 38032
rect 67660 37988 67700 37997
rect 67564 37948 67660 37988
rect 67564 37484 67604 37948
rect 67660 37920 67700 37948
rect 67755 37652 67797 37661
rect 67755 37612 67756 37652
rect 67796 37612 67797 37652
rect 67755 37603 67797 37612
rect 67756 37518 67796 37603
rect 67564 37157 67604 37444
rect 67948 37325 67988 38200
rect 68044 38191 68084 38200
rect 68140 38240 68180 38249
rect 68140 37460 68180 38200
rect 68236 38240 68276 38249
rect 68236 37661 68276 38200
rect 68332 38240 68372 38249
rect 68716 38240 68756 38249
rect 68372 38200 68564 38240
rect 68332 38191 68372 38200
rect 68235 37652 68277 37661
rect 68235 37612 68236 37652
rect 68276 37612 68277 37652
rect 68235 37603 68277 37612
rect 68140 37420 68276 37460
rect 68044 37400 68084 37409
rect 67947 37316 67989 37325
rect 67947 37276 67948 37316
rect 67988 37276 67989 37316
rect 67947 37267 67989 37276
rect 67756 37232 67796 37241
rect 67796 37192 67892 37232
rect 67756 37183 67796 37192
rect 67563 37148 67605 37157
rect 67563 37108 67564 37148
rect 67604 37108 67605 37148
rect 67563 37099 67605 37108
rect 67564 36317 67604 37099
rect 67755 36560 67797 36569
rect 67755 36520 67756 36560
rect 67796 36520 67797 36560
rect 67755 36511 67797 36520
rect 67563 36308 67605 36317
rect 67563 36268 67564 36308
rect 67604 36268 67605 36308
rect 67563 36259 67605 36268
rect 67468 36016 67604 36056
rect 67124 35848 67220 35888
rect 67276 35888 67316 35897
rect 67084 35839 67124 35848
rect 66891 35804 66933 35813
rect 66891 35764 66892 35804
rect 66932 35764 66933 35804
rect 66891 35755 66933 35764
rect 66892 35670 66932 35755
rect 66795 35384 66837 35393
rect 66795 35344 66796 35384
rect 66836 35344 66837 35384
rect 66795 35335 66837 35344
rect 66891 35300 66933 35309
rect 66891 35260 66892 35300
rect 66932 35260 66933 35300
rect 66891 35251 66933 35260
rect 66412 35216 66452 35225
rect 66603 35216 66645 35225
rect 66412 34553 66452 35176
rect 66508 35176 66604 35216
rect 66644 35176 66645 35216
rect 66411 34544 66453 34553
rect 66411 34504 66412 34544
rect 66452 34504 66453 34544
rect 66411 34495 66453 34504
rect 66219 34208 66261 34217
rect 66219 34168 66220 34208
rect 66260 34168 66261 34208
rect 66219 34159 66261 34168
rect 66220 34074 66260 34159
rect 66316 33965 66356 34336
rect 66412 34376 66452 34385
rect 66508 34376 66548 35176
rect 66603 35167 66645 35176
rect 66700 35216 66740 35225
rect 66700 34637 66740 35176
rect 66795 35216 66837 35225
rect 66795 35176 66796 35216
rect 66836 35176 66837 35216
rect 66795 35167 66837 35176
rect 66796 35082 66836 35167
rect 66699 34628 66741 34637
rect 66699 34588 66700 34628
rect 66740 34588 66741 34628
rect 66699 34579 66741 34588
rect 66452 34336 66548 34376
rect 66604 34544 66644 34553
rect 66412 34327 66452 34336
rect 66315 33956 66357 33965
rect 66315 33916 66316 33956
rect 66356 33916 66357 33956
rect 66315 33907 66357 33916
rect 66220 33704 66260 33713
rect 66604 33704 66644 34504
rect 66699 34460 66741 34469
rect 66699 34420 66700 34460
rect 66740 34420 66741 34460
rect 66699 34411 66741 34420
rect 66260 33664 66548 33704
rect 66220 33655 66260 33664
rect 66123 33620 66165 33629
rect 66123 33580 66124 33620
rect 66164 33580 66165 33620
rect 66123 33571 66165 33580
rect 66219 33536 66261 33545
rect 66219 33496 66220 33536
rect 66260 33496 66261 33536
rect 66219 33487 66261 33496
rect 66028 33412 66164 33452
rect 65164 33100 65300 33140
rect 64492 32864 64532 32873
rect 64204 32824 64492 32864
rect 64107 32276 64149 32285
rect 64107 32236 64108 32276
rect 64148 32236 64149 32276
rect 64107 32227 64149 32236
rect 64108 32213 64148 32227
rect 64108 32164 64148 32173
rect 64012 32068 64148 32108
rect 63764 31984 63956 32024
rect 63724 31975 63764 31984
rect 64011 31940 64053 31949
rect 64011 31900 64012 31940
rect 64052 31900 64053 31940
rect 64011 31891 64053 31900
rect 63628 31816 63764 31856
rect 62956 31564 63052 31604
rect 63052 31555 63092 31564
rect 63244 31564 63572 31604
rect 62764 31303 62804 31312
rect 62860 31352 62900 31361
rect 62667 31268 62709 31277
rect 62667 31228 62668 31268
rect 62708 31228 62709 31268
rect 62667 31219 62709 31228
rect 62668 31134 62708 31219
rect 62764 30848 62804 30857
rect 62860 30848 62900 31312
rect 63051 31352 63093 31361
rect 63051 31312 63052 31352
rect 63092 31312 63093 31352
rect 63051 31303 63093 31312
rect 63244 31352 63284 31564
rect 63628 31520 63668 31529
rect 63532 31480 63628 31520
rect 63357 31436 63399 31445
rect 63357 31396 63358 31436
rect 63398 31396 63399 31436
rect 63357 31387 63399 31396
rect 63244 31303 63284 31312
rect 63358 31363 63398 31387
rect 63052 31218 63092 31303
rect 63358 31301 63398 31323
rect 62804 30808 62900 30848
rect 62764 30799 62804 30808
rect 62475 30680 62517 30689
rect 62475 30640 62476 30680
rect 62516 30640 62517 30680
rect 62475 30631 62517 30640
rect 62668 30680 62708 30689
rect 62283 30596 62325 30605
rect 62283 30556 62284 30596
rect 62324 30556 62325 30596
rect 62283 30547 62325 30556
rect 62668 30428 62708 30640
rect 62859 30680 62901 30689
rect 62859 30640 62860 30680
rect 62900 30640 62901 30680
rect 62859 30631 62901 30640
rect 62956 30680 62996 30689
rect 62860 30546 62900 30631
rect 62188 30388 62708 30428
rect 61900 29791 61940 29800
rect 61707 29252 61749 29261
rect 61707 29212 61708 29252
rect 61748 29212 61749 29252
rect 61707 29203 61749 29212
rect 62668 29084 62708 30388
rect 62956 30092 62996 30640
rect 63148 30680 63188 30689
rect 63148 30428 63188 30640
rect 63532 30680 63572 31480
rect 63628 31471 63668 31480
rect 63724 30689 63764 31816
rect 64012 31806 64052 31891
rect 63532 30631 63572 30640
rect 63723 30680 63765 30689
rect 63723 30640 63724 30680
rect 63764 30640 63765 30680
rect 63723 30631 63765 30640
rect 63819 30596 63861 30605
rect 63819 30556 63820 30596
rect 63860 30556 63861 30596
rect 63819 30547 63861 30556
rect 63148 30388 63572 30428
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 63243 30092 63285 30101
rect 62956 30052 63244 30092
rect 63284 30052 63285 30092
rect 63532 30092 63572 30388
rect 63724 30092 63764 30101
rect 63532 30052 63724 30092
rect 63243 30043 63285 30052
rect 63724 30043 63764 30052
rect 63244 29840 63284 30043
rect 63339 30008 63381 30017
rect 63339 29968 63340 30008
rect 63380 29968 63381 30008
rect 63339 29959 63381 29968
rect 63340 29882 63380 29959
rect 63340 29833 63380 29842
rect 63435 29840 63477 29849
rect 63244 29791 63284 29800
rect 63435 29800 63436 29840
rect 63476 29800 63477 29840
rect 63435 29791 63477 29800
rect 63532 29840 63572 29849
rect 63724 29840 63764 29849
rect 63572 29800 63724 29840
rect 63532 29791 63572 29800
rect 63724 29791 63764 29800
rect 63436 29706 63476 29791
rect 63051 29672 63093 29681
rect 63051 29632 63052 29672
rect 63092 29632 63093 29672
rect 63051 29623 63093 29632
rect 63052 29261 63092 29623
rect 63531 29588 63573 29597
rect 63531 29548 63532 29588
rect 63572 29548 63573 29588
rect 63531 29539 63573 29548
rect 63435 29336 63477 29345
rect 63435 29296 63436 29336
rect 63476 29296 63477 29336
rect 63435 29287 63477 29296
rect 63051 29252 63093 29261
rect 63051 29212 63052 29252
rect 63092 29212 63093 29252
rect 63051 29203 63093 29212
rect 63436 29202 63476 29287
rect 63532 29168 63572 29539
rect 63820 29336 63860 30547
rect 63915 29840 63957 29849
rect 63915 29800 63916 29840
rect 63956 29800 63957 29840
rect 63915 29791 63957 29800
rect 64012 29840 64052 29849
rect 63916 29706 63956 29791
rect 64012 29345 64052 29800
rect 64011 29336 64053 29345
rect 63820 29296 63956 29336
rect 63340 29157 63380 29166
rect 63532 29119 63572 29128
rect 63628 29168 63668 29177
rect 63820 29168 63860 29177
rect 63668 29128 63820 29168
rect 63628 29119 63668 29128
rect 63340 29084 63380 29117
rect 62668 29044 63380 29084
rect 62380 29000 62420 29009
rect 61227 28412 61269 28421
rect 60940 28372 61172 28412
rect 60844 28279 60884 28288
rect 60748 28194 60788 28279
rect 61036 28160 61076 28169
rect 60843 28076 60885 28085
rect 60843 28036 60844 28076
rect 60884 28036 60885 28076
rect 60843 28027 60885 28036
rect 59692 27488 59732 27497
rect 60171 27488 60213 27497
rect 59732 27448 59924 27488
rect 59692 27439 59732 27448
rect 59500 26816 59540 26825
rect 59788 26816 59828 26825
rect 59540 26776 59636 26816
rect 59500 26767 59540 26776
rect 59308 26524 59444 26564
rect 59060 26272 59252 26312
rect 59020 26263 59060 26272
rect 58923 26144 58965 26153
rect 58923 26104 58924 26144
rect 58964 26104 58965 26144
rect 58923 26095 58965 26104
rect 59308 26121 59348 26155
rect 59404 26153 59444 26524
rect 59403 26144 59445 26153
rect 59403 26104 59404 26144
rect 59444 26104 59445 26144
rect 59403 26095 59445 26104
rect 59500 26144 59540 26153
rect 59308 26069 59348 26081
rect 58828 26011 58868 26020
rect 59307 26060 59349 26069
rect 59307 26020 59308 26060
rect 59348 26020 59349 26060
rect 59307 26011 59349 26020
rect 59211 25976 59253 25985
rect 59211 25936 59212 25976
rect 59252 25936 59253 25976
rect 59211 25927 59253 25936
rect 59020 25892 59060 25901
rect 58827 25808 58869 25817
rect 58827 25768 58828 25808
rect 58868 25768 58869 25808
rect 58827 25759 58869 25768
rect 58635 24884 58677 24893
rect 58635 24844 58636 24884
rect 58676 24844 58677 24884
rect 58635 24835 58677 24844
rect 58292 24592 58484 24632
rect 58252 24583 58292 24592
rect 58636 23876 58676 24835
rect 58732 24725 58772 25264
rect 58828 25145 58868 25759
rect 59020 25733 59060 25852
rect 59019 25724 59061 25733
rect 59019 25684 59020 25724
rect 59060 25684 59061 25724
rect 59212 25724 59252 25927
rect 59404 25892 59444 25901
rect 59500 25892 59540 26104
rect 59404 25724 59444 25852
rect 59493 25852 59540 25892
rect 59493 25808 59533 25852
rect 59493 25768 59540 25808
rect 59212 25684 59444 25724
rect 59019 25675 59061 25684
rect 59019 25556 59061 25565
rect 59019 25516 59020 25556
rect 59060 25516 59061 25556
rect 59019 25507 59061 25516
rect 58827 25136 58869 25145
rect 58827 25096 58828 25136
rect 58868 25096 58869 25136
rect 58827 25087 58869 25096
rect 58731 24716 58773 24725
rect 58731 24676 58732 24716
rect 58772 24676 58773 24716
rect 58731 24667 58773 24676
rect 58732 24548 58772 24557
rect 58828 24548 58868 25087
rect 58923 24884 58965 24893
rect 58923 24844 58924 24884
rect 58964 24844 58965 24884
rect 58923 24835 58965 24844
rect 58924 24800 58964 24835
rect 58924 24749 58964 24760
rect 58772 24508 58868 24548
rect 58732 24499 58772 24508
rect 58636 23836 58964 23876
rect 58060 23792 58100 23801
rect 58444 23792 58484 23801
rect 57964 23752 58060 23792
rect 58100 23752 58292 23792
rect 56812 23658 56852 23743
rect 57292 23658 57332 23743
rect 57676 23633 57716 23752
rect 58060 23743 58100 23752
rect 56524 23624 56564 23633
rect 56908 23624 56948 23633
rect 57388 23624 57428 23633
rect 56564 23584 56756 23624
rect 56524 23575 56564 23584
rect 56427 23288 56469 23297
rect 56427 23248 56428 23288
rect 56468 23248 56469 23288
rect 56427 23239 56469 23248
rect 56236 23020 56385 23060
rect 56044 22744 56095 22784
rect 56055 22596 56095 22744
rect 56345 22596 56385 23020
rect 56454 23036 56496 23045
rect 56454 22996 56455 23036
rect 56495 22996 56496 23036
rect 56454 22987 56496 22996
rect 56455 22596 56495 22987
rect 56716 22784 56756 23584
rect 56948 23584 57044 23624
rect 56908 23575 56948 23584
rect 56811 23288 56853 23297
rect 56811 23248 56812 23288
rect 56852 23248 56853 23288
rect 56811 23239 56853 23248
rect 56812 23060 56852 23239
rect 57004 23060 57044 23584
rect 57291 23456 57333 23465
rect 57291 23416 57292 23456
rect 57332 23416 57333 23456
rect 57291 23407 57333 23416
rect 56812 23020 56895 23060
rect 57004 23020 57185 23060
rect 56716 22744 56785 22784
rect 56745 22596 56785 22744
rect 56855 22596 56895 23020
rect 57145 22596 57185 23020
rect 57292 22784 57332 23407
rect 57388 23060 57428 23584
rect 57675 23624 57717 23633
rect 57675 23584 57676 23624
rect 57716 23584 57717 23624
rect 57675 23575 57717 23584
rect 57772 23624 57812 23633
rect 57772 23060 57812 23584
rect 58059 23624 58101 23633
rect 58059 23584 58060 23624
rect 58100 23584 58101 23624
rect 58059 23575 58101 23584
rect 58156 23624 58196 23633
rect 58060 23060 58100 23575
rect 57388 23020 57585 23060
rect 57772 23020 57985 23060
rect 57255 22744 57332 22784
rect 57255 22596 57295 22744
rect 57545 22596 57585 23020
rect 57654 22784 57696 22793
rect 57654 22744 57655 22784
rect 57695 22744 57696 22784
rect 57654 22735 57696 22744
rect 57655 22596 57695 22735
rect 57945 22596 57985 23020
rect 58055 23020 58100 23060
rect 58055 22596 58095 23020
rect 58156 22784 58196 23584
rect 58252 23060 58292 23752
rect 58444 23213 58484 23752
rect 58924 23792 58964 23836
rect 59020 23801 59060 25507
rect 59500 25304 59540 25768
rect 59596 25313 59636 26776
rect 59788 26573 59828 26776
rect 59884 26816 59924 27448
rect 60171 27448 60172 27488
rect 60212 27448 60213 27488
rect 60171 27439 60213 27448
rect 60651 27488 60693 27497
rect 60651 27448 60652 27488
rect 60692 27448 60693 27488
rect 60651 27439 60693 27448
rect 60075 27404 60117 27413
rect 60075 27364 60076 27404
rect 60116 27364 60117 27404
rect 60075 27355 60117 27364
rect 59884 26767 59924 26776
rect 59787 26564 59829 26573
rect 59787 26524 59788 26564
rect 59828 26524 59829 26564
rect 59787 26515 59829 26524
rect 59692 26144 59732 26153
rect 59116 25264 59540 25304
rect 59595 25304 59637 25313
rect 59595 25264 59596 25304
rect 59636 25264 59637 25304
rect 59116 24464 59156 25264
rect 59595 25255 59637 25264
rect 59403 25136 59445 25145
rect 59403 25096 59404 25136
rect 59444 25096 59445 25136
rect 59403 25087 59445 25096
rect 59404 24725 59444 25087
rect 59596 24893 59636 25255
rect 59595 24884 59637 24893
rect 59595 24844 59596 24884
rect 59636 24844 59637 24884
rect 59692 24884 59732 26104
rect 59788 26144 59828 26153
rect 59788 25985 59828 26104
rect 59980 26144 60020 26153
rect 60076 26144 60116 27355
rect 60172 27068 60212 27439
rect 60459 27236 60501 27245
rect 60459 27196 60460 27236
rect 60500 27196 60501 27236
rect 60459 27187 60501 27196
rect 60172 27019 60212 27028
rect 60363 26900 60405 26909
rect 60363 26860 60364 26900
rect 60404 26860 60405 26900
rect 60363 26851 60405 26860
rect 60267 26816 60309 26825
rect 60267 26776 60268 26816
rect 60308 26776 60309 26816
rect 60267 26767 60309 26776
rect 60020 26104 60212 26144
rect 59980 26095 60020 26104
rect 59787 25976 59829 25985
rect 59787 25936 59788 25976
rect 59828 25936 59829 25976
rect 59787 25927 59829 25936
rect 60172 25976 60212 26104
rect 59980 25892 60020 25901
rect 60020 25852 60116 25892
rect 59980 25843 60020 25852
rect 60076 25304 60116 25852
rect 60172 25649 60212 25936
rect 60171 25640 60213 25649
rect 60171 25600 60172 25640
rect 60212 25600 60213 25640
rect 60171 25591 60213 25600
rect 60172 25304 60212 25313
rect 60076 25264 60172 25304
rect 60172 25255 60212 25264
rect 59884 25145 59924 25230
rect 59883 25136 59925 25145
rect 59883 25096 59884 25136
rect 59924 25096 59925 25136
rect 59883 25087 59925 25096
rect 59787 24884 59829 24893
rect 59692 24844 59788 24884
rect 59828 24844 59829 24884
rect 59595 24835 59637 24844
rect 59787 24835 59829 24844
rect 60171 24884 60213 24893
rect 60171 24844 60172 24884
rect 60212 24844 60213 24884
rect 60171 24835 60213 24844
rect 59499 24800 59541 24809
rect 59499 24760 59500 24800
rect 59540 24760 59541 24800
rect 59499 24751 59541 24760
rect 59403 24716 59445 24725
rect 59403 24676 59404 24716
rect 59444 24676 59445 24716
rect 59403 24667 59445 24676
rect 59404 24582 59444 24667
rect 59500 24632 59540 24751
rect 59596 24632 59636 24835
rect 60075 24800 60117 24809
rect 60075 24760 60076 24800
rect 60116 24760 60117 24800
rect 60075 24751 60117 24760
rect 59788 24632 59828 24641
rect 59596 24592 59788 24632
rect 59500 24583 59540 24592
rect 59788 24583 59828 24592
rect 60076 24632 60116 24751
rect 60172 24716 60212 24835
rect 60172 24667 60212 24676
rect 60076 24583 60116 24592
rect 60268 24632 60308 26767
rect 60364 26766 60404 26851
rect 60460 26648 60500 27187
rect 60747 27152 60789 27161
rect 60747 27112 60748 27152
rect 60788 27112 60789 27152
rect 60747 27103 60789 27112
rect 60748 26909 60788 27103
rect 60844 27068 60884 28027
rect 60844 27019 60884 27028
rect 60940 27656 60980 27665
rect 60940 26984 60980 27616
rect 61036 27161 61076 28120
rect 61132 27245 61172 28372
rect 61227 28372 61228 28412
rect 61268 28372 61269 28412
rect 61227 28363 61269 28372
rect 61420 28412 61460 28421
rect 61228 28278 61268 28363
rect 61420 28001 61460 28372
rect 61419 27992 61461 28001
rect 61419 27952 61420 27992
rect 61460 27952 61461 27992
rect 61419 27943 61461 27952
rect 61131 27236 61173 27245
rect 61131 27196 61132 27236
rect 61172 27196 61173 27236
rect 61131 27187 61173 27196
rect 61035 27152 61077 27161
rect 61035 27112 61036 27152
rect 61076 27112 61077 27152
rect 61035 27103 61077 27112
rect 61132 26984 61172 26993
rect 60940 26944 61132 26984
rect 61132 26935 61172 26944
rect 60747 26900 60789 26909
rect 60747 26860 60748 26900
rect 60788 26860 60789 26900
rect 60747 26851 60789 26860
rect 60748 26816 60788 26851
rect 60556 26741 60596 26772
rect 60748 26766 60788 26776
rect 60940 26816 60980 26825
rect 60555 26732 60597 26741
rect 60555 26692 60556 26732
rect 60596 26692 60597 26732
rect 60555 26683 60597 26692
rect 60364 26608 60500 26648
rect 60556 26648 60596 26683
rect 60364 26237 60404 26608
rect 60556 26489 60596 26608
rect 60940 26573 60980 26776
rect 61323 26648 61365 26657
rect 61323 26608 61324 26648
rect 61364 26608 61365 26648
rect 61323 26599 61365 26608
rect 60939 26564 60981 26573
rect 60939 26524 60940 26564
rect 60980 26524 60981 26564
rect 60939 26515 60981 26524
rect 60555 26480 60597 26489
rect 60459 26440 60556 26480
rect 60596 26440 60597 26480
rect 60363 26228 60405 26237
rect 60363 26188 60364 26228
rect 60404 26188 60405 26228
rect 60363 26179 60405 26188
rect 60364 26060 60404 26179
rect 60459 26153 60499 26440
rect 60555 26431 60597 26440
rect 61131 26480 61173 26489
rect 61131 26440 61132 26480
rect 61172 26440 61173 26480
rect 61131 26431 61173 26440
rect 61132 26312 61172 26431
rect 61132 26237 61172 26272
rect 61131 26228 61173 26237
rect 61131 26188 61132 26228
rect 61172 26188 61173 26228
rect 61131 26179 61173 26188
rect 60459 26144 60501 26153
rect 60459 26104 60460 26144
rect 60500 26104 60501 26144
rect 60459 26095 60501 26104
rect 60748 26069 60788 26100
rect 60364 26011 60404 26020
rect 60555 26060 60597 26069
rect 60555 26020 60556 26060
rect 60596 26020 60597 26060
rect 60555 26011 60597 26020
rect 60747 26060 60789 26069
rect 60747 26020 60748 26060
rect 60788 26020 60789 26060
rect 60747 26011 60789 26020
rect 60940 26060 60980 26069
rect 60556 25926 60596 26011
rect 60748 25976 60788 26011
rect 60363 25892 60405 25901
rect 60363 25852 60364 25892
rect 60404 25852 60405 25892
rect 60363 25843 60405 25852
rect 60364 24800 60404 25843
rect 60748 25817 60788 25936
rect 60747 25808 60789 25817
rect 60747 25768 60748 25808
rect 60788 25768 60789 25808
rect 60747 25759 60789 25768
rect 60940 25397 60980 26020
rect 60939 25388 60981 25397
rect 60939 25348 60940 25388
rect 60980 25348 60981 25388
rect 60939 25339 60981 25348
rect 60556 25304 60596 25313
rect 60596 25264 60884 25304
rect 60556 25255 60596 25264
rect 60459 25136 60501 25145
rect 60459 25096 60460 25136
rect 60500 25096 60692 25136
rect 60459 25087 60501 25096
rect 60460 24800 60500 24809
rect 60364 24760 60460 24800
rect 60460 24751 60500 24760
rect 60268 24583 60308 24592
rect 60652 24548 60692 25096
rect 60652 24499 60692 24508
rect 59116 24415 59156 24424
rect 60844 24464 60884 25264
rect 60844 24415 60884 24424
rect 60843 23960 60885 23969
rect 60843 23920 60844 23960
rect 60884 23920 60885 23960
rect 60843 23911 60885 23920
rect 61227 23960 61269 23969
rect 61227 23920 61228 23960
rect 61268 23920 61269 23960
rect 61227 23911 61269 23920
rect 59692 23801 59732 23886
rect 60459 23876 60501 23885
rect 60459 23836 60460 23876
rect 60500 23836 60501 23876
rect 60459 23827 60501 23836
rect 60747 23876 60789 23885
rect 60747 23836 60748 23876
rect 60788 23836 60789 23876
rect 60747 23827 60789 23836
rect 58540 23624 58580 23633
rect 58443 23204 58485 23213
rect 58443 23164 58444 23204
rect 58484 23164 58485 23204
rect 58443 23155 58485 23164
rect 58540 23060 58580 23584
rect 58924 23456 58964 23752
rect 59019 23792 59061 23801
rect 59019 23752 59020 23792
rect 59060 23752 59061 23792
rect 59019 23743 59061 23752
rect 59308 23792 59348 23801
rect 59020 23624 59060 23633
rect 59060 23584 59156 23624
rect 59020 23575 59060 23584
rect 58924 23416 59060 23456
rect 58827 23204 58869 23213
rect 58827 23164 58828 23204
rect 58868 23164 58869 23204
rect 58827 23155 58869 23164
rect 58828 23060 58868 23155
rect 58252 23020 58495 23060
rect 58540 23020 58785 23060
rect 58828 23020 58895 23060
rect 58156 22744 58385 22784
rect 58345 22596 58385 22744
rect 58455 22596 58495 23020
rect 58745 22596 58785 23020
rect 58855 22596 58895 23020
rect 59020 22793 59060 23416
rect 59116 23060 59156 23584
rect 59308 23549 59348 23752
rect 59691 23792 59733 23801
rect 59691 23752 59692 23792
rect 59732 23752 59733 23792
rect 59691 23743 59733 23752
rect 59979 23792 60021 23801
rect 59979 23752 59980 23792
rect 60020 23752 60021 23792
rect 59979 23743 60021 23752
rect 60076 23792 60116 23801
rect 59404 23624 59444 23633
rect 59307 23540 59349 23549
rect 59307 23500 59308 23540
rect 59348 23500 59349 23540
rect 59307 23491 59349 23500
rect 59404 23060 59444 23584
rect 59788 23624 59828 23633
rect 59691 23540 59733 23549
rect 59691 23500 59692 23540
rect 59732 23500 59733 23540
rect 59691 23491 59733 23500
rect 59692 23060 59732 23491
rect 59116 23020 59185 23060
rect 59404 23020 59585 23060
rect 59019 22784 59061 22793
rect 59019 22744 59020 22784
rect 59060 22744 59061 22784
rect 59019 22735 59061 22744
rect 59145 22596 59185 23020
rect 59254 22784 59296 22793
rect 59254 22744 59255 22784
rect 59295 22744 59296 22784
rect 59254 22735 59296 22744
rect 59255 22596 59295 22735
rect 59545 22596 59585 23020
rect 59655 23020 59732 23060
rect 59788 23060 59828 23584
rect 59980 23060 60020 23743
rect 60076 23633 60116 23752
rect 60460 23792 60500 23827
rect 60460 23741 60500 23752
rect 60075 23624 60117 23633
rect 60075 23584 60076 23624
rect 60116 23584 60117 23624
rect 60075 23575 60117 23584
rect 60172 23624 60212 23633
rect 60172 23060 60212 23584
rect 60556 23624 60596 23633
rect 60596 23584 60692 23624
rect 60556 23575 60596 23584
rect 59788 23020 59924 23060
rect 59980 23020 60095 23060
rect 60172 23020 60308 23060
rect 59655 22596 59695 23020
rect 59884 22784 59924 23020
rect 59884 22744 59985 22784
rect 59945 22596 59985 22744
rect 60055 22596 60095 23020
rect 60268 22784 60308 23020
rect 60652 22868 60692 23584
rect 60748 23060 60788 23827
rect 60844 23792 60884 23911
rect 60844 23743 60884 23752
rect 60940 23624 60980 23633
rect 60940 23060 60980 23584
rect 61228 23060 61268 23911
rect 61324 23792 61364 26599
rect 61419 26144 61461 26153
rect 61419 26104 61420 26144
rect 61460 26104 61461 26144
rect 61419 26095 61461 26104
rect 61420 25304 61460 26095
rect 61516 25901 61556 28531
rect 61612 28421 61652 28540
rect 62284 28960 62380 29000
rect 61611 28412 61653 28421
rect 61611 28372 61612 28412
rect 61652 28372 61653 28412
rect 61611 28363 61653 28372
rect 61803 28328 61845 28337
rect 61803 28288 61804 28328
rect 61844 28288 61845 28328
rect 61803 28279 61845 28288
rect 62284 28328 62324 28960
rect 62380 28951 62420 28960
rect 62284 28279 62324 28288
rect 61804 27656 61844 28279
rect 61900 28244 61940 28253
rect 61900 27833 61940 28204
rect 61899 27824 61941 27833
rect 61899 27784 61900 27824
rect 61940 27784 61941 27824
rect 61899 27775 61941 27784
rect 61611 26648 61653 26657
rect 61611 26608 61612 26648
rect 61652 26608 61653 26648
rect 61611 26599 61653 26608
rect 61612 26489 61652 26599
rect 61611 26480 61653 26489
rect 61611 26440 61612 26480
rect 61652 26440 61653 26480
rect 61611 26431 61653 26440
rect 61611 26228 61653 26237
rect 61611 26188 61612 26228
rect 61652 26188 61653 26228
rect 61611 26179 61653 26188
rect 61612 26094 61652 26179
rect 61804 26153 61844 27616
rect 61899 27068 61941 27077
rect 61899 27028 61900 27068
rect 61940 27028 61941 27068
rect 61899 27019 61941 27028
rect 61900 26825 61940 27019
rect 62092 26984 62132 26993
rect 61899 26816 61941 26825
rect 61899 26776 61900 26816
rect 61940 26776 61941 26816
rect 61899 26767 61941 26776
rect 61803 26144 61845 26153
rect 61803 26104 61804 26144
rect 61844 26104 61845 26144
rect 61803 26095 61845 26104
rect 61996 26144 62036 26153
rect 62092 26144 62132 26944
rect 62860 26825 62900 29044
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 63147 28328 63189 28337
rect 63147 28288 63148 28328
rect 63188 28288 63189 28328
rect 63147 28279 63189 28288
rect 63148 28194 63188 28279
rect 63820 28253 63860 29128
rect 63916 29168 63956 29296
rect 64011 29296 64012 29336
rect 64052 29296 64053 29336
rect 64108 29336 64148 32068
rect 64204 31697 64244 32824
rect 64492 32815 64532 32824
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 64491 32360 64533 32369
rect 64491 32320 64492 32360
rect 64532 32320 64533 32360
rect 64491 32311 64533 32320
rect 64300 32192 64340 32201
rect 64300 32033 64340 32152
rect 64492 32192 64532 32311
rect 64779 32276 64821 32285
rect 64779 32236 64780 32276
rect 64820 32236 64821 32276
rect 64779 32227 64821 32236
rect 64492 32143 64532 32152
rect 64299 32024 64341 32033
rect 64299 31984 64300 32024
rect 64340 31984 64341 32024
rect 64299 31975 64341 31984
rect 64396 31940 64436 31949
rect 64203 31688 64245 31697
rect 64203 31648 64204 31688
rect 64244 31648 64245 31688
rect 64203 31639 64245 31648
rect 64396 31445 64436 31900
rect 64395 31436 64437 31445
rect 64395 31396 64396 31436
rect 64436 31396 64437 31436
rect 64395 31387 64437 31396
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 64780 30848 64820 32227
rect 65163 31940 65205 31949
rect 65163 31900 65164 31940
rect 65204 31900 65205 31940
rect 65163 31891 65205 31900
rect 64684 30808 64820 30848
rect 64395 30680 64437 30689
rect 64395 30640 64396 30680
rect 64436 30640 64437 30680
rect 64395 30631 64437 30640
rect 64203 30596 64245 30605
rect 64203 30556 64204 30596
rect 64244 30556 64245 30596
rect 64203 30547 64245 30556
rect 64204 29513 64244 30547
rect 64396 30546 64436 30631
rect 64684 29840 64724 30808
rect 65068 30008 65108 30017
rect 64780 29849 64820 29880
rect 64684 29791 64724 29800
rect 64779 29840 64821 29849
rect 64779 29800 64780 29840
rect 64820 29800 64821 29840
rect 64779 29791 64821 29800
rect 64876 29840 64916 29849
rect 65068 29840 65108 29968
rect 64916 29800 65108 29840
rect 64876 29791 64916 29800
rect 64780 29756 64820 29791
rect 64203 29504 64245 29513
rect 64203 29464 64204 29504
rect 64244 29464 64245 29504
rect 64203 29455 64245 29464
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 64108 29296 64244 29336
rect 64011 29287 64053 29296
rect 64204 29177 64244 29296
rect 64780 29177 64820 29716
rect 63819 28244 63861 28253
rect 63819 28204 63820 28244
rect 63860 28204 63861 28244
rect 63819 28195 63861 28204
rect 63916 27992 63956 29128
rect 64011 29168 64053 29177
rect 64011 29128 64012 29168
rect 64052 29128 64053 29168
rect 64011 29119 64053 29128
rect 64108 29168 64148 29177
rect 64012 29034 64052 29119
rect 63628 27952 63956 27992
rect 62956 27404 62996 27413
rect 62859 26816 62901 26825
rect 62859 26776 62860 26816
rect 62900 26776 62901 26816
rect 62859 26767 62901 26776
rect 62956 26573 62996 27364
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 63628 26993 63668 27952
rect 63915 27824 63957 27833
rect 63915 27784 63916 27824
rect 63956 27784 63957 27824
rect 63915 27775 63957 27784
rect 63916 27690 63956 27775
rect 63724 27656 63764 27665
rect 63724 27068 63764 27616
rect 63819 27656 63861 27665
rect 63819 27616 63820 27656
rect 63860 27616 63861 27656
rect 63819 27607 63861 27616
rect 64012 27656 64052 27665
rect 64108 27656 64148 29128
rect 64203 29168 64245 29177
rect 64203 29128 64204 29168
rect 64244 29128 64245 29168
rect 64203 29119 64245 29128
rect 64779 29168 64821 29177
rect 64779 29128 64780 29168
rect 64820 29128 64821 29168
rect 64779 29119 64821 29128
rect 65067 28832 65109 28841
rect 65067 28792 65068 28832
rect 65108 28792 65109 28832
rect 65067 28783 65109 28792
rect 64492 28496 64532 28505
rect 64532 28456 64724 28496
rect 64492 28447 64532 28456
rect 64299 28244 64341 28253
rect 64299 28204 64300 28244
rect 64340 28204 64341 28244
rect 64299 28195 64341 28204
rect 64300 28160 64340 28195
rect 64684 28160 64724 28456
rect 64780 28337 64820 28422
rect 64779 28328 64821 28337
rect 64779 28288 64780 28328
rect 64820 28288 64821 28328
rect 64779 28279 64821 28288
rect 64876 28328 64916 28337
rect 65068 28328 65108 28783
rect 65164 28505 65204 31891
rect 65163 28496 65205 28505
rect 65163 28456 65164 28496
rect 65204 28456 65205 28496
rect 65260 28496 65300 33100
rect 66027 32864 66069 32873
rect 66027 32824 66028 32864
rect 66068 32824 66069 32864
rect 66027 32815 66069 32824
rect 66124 32864 66164 33412
rect 66124 32815 66164 32824
rect 66220 32864 66260 33487
rect 66508 33116 66548 33664
rect 66604 33655 66644 33664
rect 66700 33140 66740 34411
rect 66795 34208 66837 34217
rect 66795 34168 66796 34208
rect 66836 34168 66837 34208
rect 66795 34159 66837 34168
rect 66508 33067 66548 33076
rect 66604 33100 66740 33140
rect 66220 32815 66260 32824
rect 66316 32864 66356 32873
rect 66508 32864 66548 32873
rect 66356 32824 66508 32864
rect 66316 32815 66356 32824
rect 66508 32815 66548 32824
rect 65643 32696 65685 32705
rect 65643 32656 65644 32696
rect 65684 32656 65685 32696
rect 65643 32647 65685 32656
rect 65355 32528 65397 32537
rect 65355 32488 65356 32528
rect 65396 32488 65397 32528
rect 65355 32479 65397 32488
rect 65356 32285 65396 32479
rect 65644 32369 65684 32647
rect 65931 32612 65973 32621
rect 65931 32572 65932 32612
rect 65972 32572 65973 32612
rect 65931 32563 65973 32572
rect 65643 32360 65685 32369
rect 65643 32320 65644 32360
rect 65684 32320 65685 32360
rect 65643 32311 65685 32320
rect 65355 32276 65397 32285
rect 65355 32236 65356 32276
rect 65396 32236 65397 32276
rect 65355 32227 65397 32236
rect 65356 32192 65396 32227
rect 65356 32142 65396 32152
rect 65548 32192 65588 32201
rect 65588 32152 65780 32192
rect 65548 32143 65588 32152
rect 65451 32024 65493 32033
rect 65451 31984 65452 32024
rect 65492 31984 65493 32024
rect 65451 31975 65493 31984
rect 65740 32024 65780 32152
rect 65740 31975 65780 31984
rect 65452 31890 65492 31975
rect 65932 30848 65972 32563
rect 66028 32276 66068 32815
rect 66604 32696 66644 33100
rect 66412 32656 66644 32696
rect 66700 32864 66740 32873
rect 66219 32444 66261 32453
rect 66219 32404 66220 32444
rect 66260 32404 66261 32444
rect 66219 32395 66261 32404
rect 66028 32227 66068 32236
rect 66124 32192 66164 32201
rect 66124 31949 66164 32152
rect 66123 31940 66165 31949
rect 66123 31900 66124 31940
rect 66164 31900 66165 31940
rect 66123 31891 66165 31900
rect 65932 30808 66068 30848
rect 65835 30764 65877 30773
rect 65835 30724 65836 30764
rect 65876 30724 65877 30764
rect 65835 30715 65877 30724
rect 65548 30428 65588 30437
rect 65548 30269 65588 30388
rect 65355 30260 65397 30269
rect 65355 30220 65356 30260
rect 65396 30220 65397 30260
rect 65355 30211 65397 30220
rect 65547 30260 65589 30269
rect 65547 30220 65548 30260
rect 65588 30220 65589 30260
rect 65547 30211 65589 30220
rect 65356 29840 65396 30211
rect 65836 29849 65876 30715
rect 65932 30680 65972 30691
rect 65932 30605 65972 30640
rect 65931 30596 65973 30605
rect 65931 30556 65932 30596
rect 65972 30556 65973 30596
rect 66028 30596 66068 30808
rect 66124 30773 66164 30788
rect 66123 30764 66165 30773
rect 66123 30724 66124 30764
rect 66164 30724 66165 30764
rect 66123 30715 66165 30724
rect 66124 30693 66164 30715
rect 66124 30644 66164 30653
rect 66028 30556 66164 30596
rect 65931 30547 65973 30556
rect 66028 30428 66068 30437
rect 65932 30388 66028 30428
rect 65356 29791 65396 29800
rect 65451 29840 65493 29849
rect 65740 29840 65780 29849
rect 65451 29800 65452 29840
rect 65492 29800 65493 29840
rect 65451 29791 65493 29800
rect 65548 29800 65740 29840
rect 65452 29706 65492 29791
rect 65548 28841 65588 29800
rect 65740 29791 65780 29800
rect 65835 29840 65877 29849
rect 65835 29800 65836 29840
rect 65876 29800 65877 29840
rect 65835 29791 65877 29800
rect 65643 29336 65685 29345
rect 65643 29296 65644 29336
rect 65684 29296 65685 29336
rect 65643 29287 65685 29296
rect 65644 29168 65684 29287
rect 65547 28832 65589 28841
rect 65547 28792 65548 28832
rect 65588 28792 65589 28832
rect 65547 28783 65589 28792
rect 65260 28456 65588 28496
rect 65163 28447 65205 28456
rect 65164 28328 65204 28337
rect 65068 28288 65164 28328
rect 64684 28120 64785 28160
rect 64300 28109 64340 28120
rect 64745 28076 64785 28120
rect 64745 28036 64820 28076
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 64052 27616 64148 27656
rect 64780 27656 64820 28036
rect 64876 27833 64916 28288
rect 65164 28279 65204 28288
rect 65259 28160 65301 28169
rect 65259 28120 65260 28160
rect 65300 28120 65301 28160
rect 65259 28111 65301 28120
rect 65067 28076 65109 28085
rect 65067 28036 65068 28076
rect 65108 28036 65109 28076
rect 65067 28027 65109 28036
rect 64875 27824 64917 27833
rect 64875 27784 64876 27824
rect 64916 27784 64917 27824
rect 64875 27775 64917 27784
rect 64012 27607 64052 27616
rect 64780 27607 64820 27616
rect 64875 27656 64917 27665
rect 64875 27616 64876 27656
rect 64916 27616 64917 27656
rect 64875 27607 64917 27616
rect 64972 27656 65012 27665
rect 63820 27522 63860 27607
rect 64876 27522 64916 27607
rect 63820 27068 63860 27077
rect 63724 27028 63820 27068
rect 63820 27019 63860 27028
rect 63627 26984 63669 26993
rect 63627 26944 63628 26984
rect 63668 26944 63669 26984
rect 63627 26935 63669 26944
rect 64203 26984 64245 26993
rect 64203 26944 64204 26984
rect 64244 26944 64245 26984
rect 64012 26909 64052 26940
rect 64203 26935 64245 26944
rect 64011 26900 64053 26909
rect 64011 26860 64012 26900
rect 64052 26860 64053 26900
rect 64011 26851 64053 26860
rect 63819 26816 63861 26825
rect 63819 26776 63820 26816
rect 63860 26776 63861 26816
rect 63819 26767 63861 26776
rect 64012 26816 64052 26851
rect 62955 26564 62997 26573
rect 62955 26524 62956 26564
rect 62996 26524 62997 26564
rect 62955 26515 62997 26524
rect 63531 26312 63573 26321
rect 63531 26272 63532 26312
rect 63572 26272 63573 26312
rect 63531 26263 63573 26272
rect 62036 26104 62132 26144
rect 62859 26144 62901 26153
rect 62859 26104 62860 26144
rect 62900 26104 62901 26144
rect 61996 26095 62036 26104
rect 62859 26095 62901 26104
rect 62860 26010 62900 26095
rect 61515 25892 61557 25901
rect 61515 25852 61516 25892
rect 61556 25852 61557 25892
rect 61515 25843 61557 25852
rect 61420 25255 61460 25264
rect 61516 25145 61556 25843
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 63532 25556 63572 26263
rect 63820 26153 63860 26767
rect 64012 26573 64052 26776
rect 64108 26816 64148 26825
rect 64011 26564 64053 26573
rect 64011 26524 64012 26564
rect 64052 26524 64053 26564
rect 64011 26515 64053 26524
rect 63819 26144 63861 26153
rect 63819 26104 63820 26144
rect 63860 26104 63861 26144
rect 63819 26095 63861 26104
rect 64012 25892 64052 25901
rect 64108 25892 64148 26776
rect 64204 26312 64244 26935
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 64395 26312 64437 26321
rect 64204 26272 64340 26312
rect 64204 26144 64244 26153
rect 64204 25892 64244 26104
rect 64300 26144 64340 26272
rect 64395 26272 64396 26312
rect 64436 26272 64437 26312
rect 64972 26312 65012 27616
rect 65068 27488 65108 28027
rect 65163 27992 65205 28001
rect 65163 27952 65164 27992
rect 65204 27952 65205 27992
rect 65163 27943 65205 27952
rect 65164 27656 65204 27943
rect 65164 27607 65204 27616
rect 65164 27488 65204 27497
rect 65068 27448 65164 27488
rect 65164 27439 65204 27448
rect 65260 27413 65300 28111
rect 65355 27656 65397 27665
rect 65355 27616 65356 27656
rect 65396 27616 65397 27656
rect 65355 27607 65397 27616
rect 65452 27656 65492 27667
rect 65356 27522 65396 27607
rect 65452 27581 65492 27616
rect 65451 27572 65493 27581
rect 65451 27532 65452 27572
rect 65492 27532 65493 27572
rect 65451 27523 65493 27532
rect 65259 27404 65301 27413
rect 65259 27364 65260 27404
rect 65300 27364 65301 27404
rect 65259 27355 65301 27364
rect 65163 27320 65205 27329
rect 65163 27280 65164 27320
rect 65204 27280 65205 27320
rect 65163 27271 65205 27280
rect 64972 26272 65108 26312
rect 64395 26263 64437 26272
rect 64300 26095 64340 26104
rect 64396 26144 64436 26263
rect 64779 26228 64821 26237
rect 64779 26188 64780 26228
rect 64820 26188 64821 26228
rect 64779 26179 64821 26188
rect 64396 26095 64436 26104
rect 64492 26144 64532 26153
rect 64684 26144 64724 26153
rect 64532 26104 64684 26144
rect 64492 26095 64532 26104
rect 64684 26095 64724 26104
rect 64780 26094 64820 26179
rect 64876 26144 64916 26153
rect 64299 25976 64341 25985
rect 64299 25936 64300 25976
rect 64340 25936 64341 25976
rect 64299 25927 64341 25936
rect 64779 25976 64821 25985
rect 64876 25976 64916 26104
rect 64972 26144 65012 26153
rect 64972 25985 65012 26104
rect 64779 25936 64780 25976
rect 64820 25936 64916 25976
rect 64971 25976 65013 25985
rect 64971 25936 64972 25976
rect 65012 25936 65013 25976
rect 64779 25927 64821 25936
rect 64971 25927 65013 25936
rect 64052 25852 64244 25892
rect 64012 25808 64052 25852
rect 63436 25516 63572 25556
rect 63724 25768 64052 25808
rect 63436 25472 63476 25516
rect 63244 25432 63476 25472
rect 63147 25304 63189 25313
rect 63147 25264 63148 25304
rect 63188 25264 63189 25304
rect 63147 25255 63189 25264
rect 63148 25170 63188 25255
rect 61515 25136 61557 25145
rect 61515 25096 61516 25136
rect 61556 25096 61557 25136
rect 61515 25087 61557 25096
rect 62572 25136 62612 25145
rect 61707 25052 61749 25061
rect 61707 25012 61708 25052
rect 61748 25012 61749 25052
rect 61707 25003 61749 25012
rect 61708 23792 61748 25003
rect 62572 24809 62612 25096
rect 62571 24800 62613 24809
rect 62571 24760 62572 24800
rect 62612 24760 62613 24800
rect 62571 24751 62613 24760
rect 62475 24296 62517 24305
rect 62475 24256 62476 24296
rect 62516 24256 62517 24296
rect 62475 24247 62517 24256
rect 62091 24044 62133 24053
rect 62091 24004 62092 24044
rect 62132 24004 62133 24044
rect 62091 23995 62133 24004
rect 62092 23792 62132 23995
rect 62476 23792 62516 24247
rect 62572 24053 62612 24751
rect 62571 24044 62613 24053
rect 62571 24004 62572 24044
rect 62612 24004 62613 24044
rect 62571 23995 62613 24004
rect 63244 23969 63284 25432
rect 63435 25304 63477 25313
rect 63435 25264 63436 25304
rect 63476 25264 63477 25304
rect 63435 25255 63477 25264
rect 63532 25304 63572 25313
rect 63724 25304 63764 25768
rect 63572 25264 63764 25304
rect 63820 25472 63860 25481
rect 63532 25255 63572 25264
rect 63436 25170 63476 25255
rect 63531 25136 63573 25145
rect 63531 25096 63532 25136
rect 63572 25096 63573 25136
rect 63531 25087 63573 25096
rect 63435 24968 63477 24977
rect 63435 24928 63436 24968
rect 63476 24928 63477 24968
rect 63435 24919 63477 24928
rect 63243 23960 63285 23969
rect 63243 23920 63244 23960
rect 63284 23920 63285 23960
rect 63436 23960 63476 24919
rect 63532 24632 63572 25087
rect 63532 24583 63572 24592
rect 63627 24632 63669 24641
rect 63627 24592 63628 24632
rect 63668 24592 63669 24632
rect 63627 24583 63669 24592
rect 63724 24632 63764 24641
rect 63820 24632 63860 25432
rect 63915 25304 63957 25313
rect 63915 25264 63916 25304
rect 63956 25264 63957 25304
rect 63915 25255 63957 25264
rect 63916 24893 63956 25255
rect 64012 25220 64052 25229
rect 63915 24884 63957 24893
rect 63915 24844 63916 24884
rect 63956 24844 63957 24884
rect 63915 24835 63957 24844
rect 64012 24800 64052 25180
rect 64300 25136 64340 25927
rect 65068 25733 65108 26272
rect 65067 25724 65109 25733
rect 65067 25684 65068 25724
rect 65108 25684 65109 25724
rect 65067 25675 65109 25684
rect 64396 25304 64436 25313
rect 64436 25264 64820 25304
rect 64396 25255 64436 25264
rect 64012 24751 64052 24760
rect 64108 25096 64340 25136
rect 63915 24716 63957 24725
rect 63915 24676 63916 24716
rect 63956 24676 63957 24716
rect 63915 24667 63957 24676
rect 63764 24592 63860 24632
rect 63916 24632 63956 24667
rect 64108 24641 64148 25096
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 64204 24760 64532 24800
rect 63724 24583 63764 24592
rect 63628 24498 63668 24583
rect 63916 24581 63956 24592
rect 64107 24632 64149 24641
rect 64107 24592 64108 24632
rect 64148 24592 64149 24632
rect 64107 24583 64149 24592
rect 64204 24632 64244 24760
rect 64492 24716 64532 24760
rect 64492 24667 64532 24676
rect 64587 24716 64629 24725
rect 64587 24676 64588 24716
rect 64628 24676 64629 24716
rect 64587 24667 64629 24676
rect 64204 24583 64244 24592
rect 64395 24632 64437 24641
rect 64395 24592 64396 24632
rect 64436 24592 64437 24632
rect 64395 24583 64437 24592
rect 64588 24632 64628 24667
rect 64108 24498 64148 24583
rect 64396 24498 64436 24583
rect 64588 24581 64628 24592
rect 64491 24464 64533 24473
rect 64491 24424 64492 24464
rect 64532 24424 64533 24464
rect 64491 24415 64533 24424
rect 64780 24464 64820 25264
rect 65068 25145 65108 25675
rect 65067 25136 65109 25145
rect 65067 25096 65068 25136
rect 65108 25096 65109 25136
rect 65067 25087 65109 25096
rect 65164 24968 65204 27271
rect 65260 25304 65300 27355
rect 65548 26816 65588 28456
rect 65644 28001 65684 29128
rect 65740 29252 65780 29261
rect 65740 29000 65780 29212
rect 65836 29177 65876 29262
rect 65835 29168 65877 29177
rect 65835 29128 65836 29168
rect 65876 29128 65877 29168
rect 65835 29119 65877 29128
rect 65932 29168 65972 30388
rect 66028 30379 66068 30388
rect 65932 29119 65972 29128
rect 66028 29756 66068 29765
rect 66028 29000 66068 29716
rect 65740 28960 66068 29000
rect 66124 28580 66164 30556
rect 65932 28540 66164 28580
rect 65740 28244 65780 28253
rect 65740 28085 65780 28204
rect 65739 28076 65781 28085
rect 65739 28036 65740 28076
rect 65780 28036 65781 28076
rect 65739 28027 65781 28036
rect 65932 28001 65972 28540
rect 66220 28496 66260 32395
rect 66412 32192 66452 32656
rect 66700 32360 66740 32824
rect 66796 32864 66836 34159
rect 66796 32815 66836 32824
rect 66892 32537 66932 35251
rect 66988 34880 67028 35839
rect 67276 35309 67316 35848
rect 67371 35888 67413 35897
rect 67371 35848 67372 35888
rect 67412 35848 67413 35888
rect 67371 35839 67413 35848
rect 67468 35888 67508 35897
rect 67372 35754 67412 35839
rect 67468 35468 67508 35848
rect 67372 35428 67508 35468
rect 67275 35300 67317 35309
rect 67275 35260 67276 35300
rect 67316 35260 67317 35300
rect 67275 35251 67317 35260
rect 67084 35048 67124 35057
rect 67372 35048 67412 35428
rect 67124 35008 67412 35048
rect 67468 35216 67508 35225
rect 67084 34999 67124 35008
rect 66988 34840 67124 34880
rect 66987 34712 67029 34721
rect 66987 34672 66988 34712
rect 67028 34672 67029 34712
rect 66987 34663 67029 34672
rect 66988 34628 67028 34663
rect 66988 34577 67028 34588
rect 66988 34376 67028 34385
rect 67084 34376 67124 34840
rect 67468 34721 67508 35176
rect 67467 34712 67509 34721
rect 67467 34672 67468 34712
rect 67508 34672 67509 34712
rect 67467 34663 67509 34672
rect 67564 34544 67604 36016
rect 67659 34628 67701 34637
rect 67659 34588 67660 34628
rect 67700 34588 67701 34628
rect 67659 34579 67701 34588
rect 67372 34504 67604 34544
rect 67180 34376 67220 34385
rect 67084 34336 67180 34376
rect 66891 32528 66933 32537
rect 66891 32488 66892 32528
rect 66932 32488 66933 32528
rect 66891 32479 66933 32488
rect 66891 32360 66933 32369
rect 66700 32320 66836 32360
rect 66700 32192 66740 32201
rect 66316 32152 66412 32192
rect 66316 28841 66356 32152
rect 66412 32143 66452 32152
rect 66508 32152 66700 32192
rect 66412 31604 66452 31613
rect 66508 31604 66548 32152
rect 66700 32143 66740 32152
rect 66603 32024 66645 32033
rect 66796 32024 66836 32320
rect 66891 32320 66892 32360
rect 66932 32320 66933 32360
rect 66891 32311 66933 32320
rect 66603 31984 66604 32024
rect 66644 31984 66836 32024
rect 66603 31975 66645 31984
rect 66452 31564 66548 31604
rect 66412 31555 66452 31564
rect 66411 31436 66453 31445
rect 66411 31396 66412 31436
rect 66452 31396 66453 31436
rect 66411 31387 66453 31396
rect 66412 31352 66452 31387
rect 66412 31301 66452 31312
rect 66604 31352 66644 31975
rect 66795 31436 66837 31445
rect 66795 31396 66796 31436
rect 66836 31396 66837 31436
rect 66795 31387 66837 31396
rect 66604 31303 66644 31312
rect 66700 31352 66740 31363
rect 66700 31277 66740 31312
rect 66699 31268 66741 31277
rect 66699 31228 66700 31268
rect 66740 31228 66741 31268
rect 66699 31219 66741 31228
rect 66603 31100 66645 31109
rect 66603 31060 66604 31100
rect 66644 31060 66645 31100
rect 66603 31051 66645 31060
rect 66508 30512 66548 30521
rect 66412 30472 66508 30512
rect 66412 29840 66452 30472
rect 66508 30463 66548 30472
rect 66412 29791 66452 29800
rect 66315 28832 66357 28841
rect 66315 28792 66316 28832
rect 66356 28792 66357 28832
rect 66315 28783 66357 28792
rect 66028 28456 66260 28496
rect 65643 27992 65685 28001
rect 65643 27952 65644 27992
rect 65684 27952 65685 27992
rect 65643 27943 65685 27952
rect 65931 27992 65973 28001
rect 65931 27952 65932 27992
rect 65972 27952 65973 27992
rect 65931 27943 65973 27952
rect 65644 27784 65972 27824
rect 65644 27656 65684 27784
rect 65644 27607 65684 27616
rect 65835 27656 65877 27665
rect 65835 27616 65836 27656
rect 65876 27616 65877 27656
rect 65835 27607 65877 27616
rect 65739 27572 65781 27581
rect 65739 27532 65740 27572
rect 65780 27532 65781 27572
rect 65739 27523 65781 27532
rect 65740 27438 65780 27523
rect 65836 27522 65876 27607
rect 65548 26776 65780 26816
rect 65644 26648 65684 26657
rect 65547 26564 65589 26573
rect 65547 26524 65548 26564
rect 65588 26524 65589 26564
rect 65547 26515 65589 26524
rect 65356 26153 65396 26238
rect 65355 26144 65397 26153
rect 65355 26104 65356 26144
rect 65396 26104 65397 26144
rect 65355 26095 65397 26104
rect 65548 26144 65588 26515
rect 65644 26153 65684 26608
rect 65355 25976 65397 25985
rect 65355 25936 65356 25976
rect 65396 25936 65397 25976
rect 65355 25927 65397 25936
rect 65356 25842 65396 25927
rect 65260 25255 65300 25264
rect 64780 24415 64820 24424
rect 64876 24928 65204 24968
rect 63436 23920 63764 23960
rect 63243 23911 63285 23920
rect 62860 23792 62900 23801
rect 61364 23752 61652 23792
rect 61324 23743 61364 23752
rect 61420 23624 61460 23633
rect 61420 23060 61460 23584
rect 61612 23060 61652 23752
rect 61748 23752 62036 23792
rect 61708 23743 61748 23752
rect 61804 23624 61844 23633
rect 61804 23060 61844 23584
rect 61996 23060 62036 23752
rect 62132 23752 62420 23792
rect 62092 23743 62132 23752
rect 62188 23624 62228 23633
rect 62188 23060 62228 23584
rect 62380 23060 62420 23752
rect 62476 23633 62516 23752
rect 62764 23752 62860 23792
rect 62475 23624 62517 23633
rect 62475 23584 62476 23624
rect 62516 23584 62517 23624
rect 62475 23575 62517 23584
rect 62572 23624 62612 23633
rect 62572 23060 62612 23584
rect 62764 23381 62804 23752
rect 62860 23743 62900 23752
rect 63244 23792 63284 23803
rect 63244 23717 63284 23752
rect 63724 23792 63764 23920
rect 64107 23792 64149 23801
rect 64492 23792 64532 24415
rect 64876 23792 64916 24928
rect 65548 24641 65588 26104
rect 65643 26144 65685 26153
rect 65643 26104 65644 26144
rect 65684 26104 65685 26144
rect 65643 26095 65685 26104
rect 65644 26010 65684 26095
rect 65547 24632 65589 24641
rect 65547 24592 65548 24632
rect 65588 24592 65589 24632
rect 65547 24583 65589 24592
rect 65259 23960 65301 23969
rect 65259 23920 65260 23960
rect 65300 23920 65301 23960
rect 65259 23911 65301 23920
rect 65643 23960 65685 23969
rect 65643 23920 65644 23960
rect 65684 23920 65685 23960
rect 65643 23911 65685 23920
rect 65260 23792 65300 23911
rect 63764 23752 64052 23792
rect 63724 23743 63764 23752
rect 63243 23708 63285 23717
rect 63243 23668 63244 23708
rect 63284 23668 63285 23708
rect 63243 23659 63285 23668
rect 63627 23708 63669 23717
rect 63627 23668 63628 23708
rect 63668 23668 63669 23708
rect 63627 23659 63669 23668
rect 62859 23624 62901 23633
rect 62859 23584 62860 23624
rect 62900 23584 62901 23624
rect 62859 23575 62901 23584
rect 62956 23624 62996 23633
rect 62763 23372 62805 23381
rect 62763 23332 62764 23372
rect 62804 23332 62805 23372
rect 62763 23323 62805 23332
rect 62860 23060 62900 23575
rect 60748 23020 60895 23060
rect 60940 23020 61185 23060
rect 61228 23020 61295 23060
rect 61420 23020 61556 23060
rect 61612 23020 61695 23060
rect 61804 23020 61940 23060
rect 61996 23020 62095 23060
rect 62188 23020 62324 23060
rect 62380 23020 62495 23060
rect 62572 23020 62785 23060
rect 60652 22828 60785 22868
rect 60464 22793 60504 22815
rect 60463 22784 60505 22793
rect 60268 22744 60385 22784
rect 60345 22596 60385 22744
rect 60455 22744 60464 22784
rect 60504 22744 60505 22784
rect 60455 22735 60505 22744
rect 60455 22596 60495 22735
rect 60745 22596 60785 22828
rect 60855 22596 60895 23020
rect 61145 22596 61185 23020
rect 61255 22596 61295 23020
rect 61516 22784 61556 23020
rect 61516 22744 61585 22784
rect 61545 22596 61585 22744
rect 61655 22596 61695 23020
rect 61900 22784 61940 23020
rect 61900 22744 61985 22784
rect 61945 22596 61985 22744
rect 62055 22596 62095 23020
rect 62284 22784 62324 23020
rect 62284 22744 62385 22784
rect 62345 22596 62385 22744
rect 62455 22596 62495 23020
rect 62745 22596 62785 23020
rect 62855 23020 62900 23060
rect 62956 23060 62996 23584
rect 63340 23624 63380 23633
rect 63380 23584 63476 23624
rect 63340 23575 63380 23584
rect 63243 23372 63285 23381
rect 63243 23332 63244 23372
rect 63284 23332 63285 23372
rect 63243 23323 63285 23332
rect 63244 23060 63284 23323
rect 63436 23060 63476 23584
rect 63628 23060 63668 23659
rect 63820 23624 63860 23633
rect 63820 23060 63860 23584
rect 64012 23060 64052 23752
rect 64107 23752 64108 23792
rect 64148 23752 64436 23792
rect 64107 23743 64149 23752
rect 64108 23658 64148 23743
rect 64204 23624 64244 23633
rect 64204 23060 64244 23584
rect 64396 23060 64436 23752
rect 64532 23752 64820 23792
rect 64492 23743 64532 23752
rect 64588 23624 64628 23633
rect 64588 23060 64628 23584
rect 64780 23060 64820 23752
rect 64916 23752 65204 23792
rect 64876 23743 64916 23752
rect 64972 23624 65012 23633
rect 64972 23060 65012 23584
rect 65164 23540 65204 23752
rect 65260 23743 65300 23752
rect 65356 23624 65396 23633
rect 65164 23500 65300 23540
rect 65260 23060 65300 23500
rect 62956 23020 63185 23060
rect 63244 23020 63295 23060
rect 63436 23020 63585 23060
rect 63628 23020 63695 23060
rect 63820 23020 63956 23060
rect 64012 23020 64095 23060
rect 64204 23020 64340 23060
rect 64396 23020 64495 23060
rect 64588 23020 64724 23060
rect 64780 23020 64895 23060
rect 64972 23020 65185 23060
rect 62855 22596 62895 23020
rect 63145 22596 63185 23020
rect 63255 22596 63295 23020
rect 63545 22596 63585 23020
rect 63655 22596 63695 23020
rect 63916 22784 63956 23020
rect 63916 22744 63985 22784
rect 63945 22596 63985 22744
rect 64055 22596 64095 23020
rect 64300 22784 64340 23020
rect 64300 22744 64385 22784
rect 64345 22596 64385 22744
rect 64455 22596 64495 23020
rect 64684 22784 64724 23020
rect 64684 22744 64785 22784
rect 64745 22596 64785 22744
rect 64855 22596 64895 23020
rect 65145 22596 65185 23020
rect 65255 23020 65300 23060
rect 65356 23060 65396 23584
rect 65644 23060 65684 23911
rect 65740 23792 65780 26776
rect 65932 26573 65972 27784
rect 65931 26564 65973 26573
rect 65931 26524 65932 26564
rect 65972 26524 65973 26564
rect 65931 26515 65973 26524
rect 66028 23969 66068 28456
rect 66124 28328 66164 28337
rect 66164 28288 66260 28328
rect 66124 28279 66164 28288
rect 66123 27992 66165 28001
rect 66123 27952 66124 27992
rect 66164 27952 66165 27992
rect 66123 27943 66165 27952
rect 66027 23960 66069 23969
rect 66027 23920 66028 23960
rect 66068 23920 66069 23960
rect 66027 23911 66069 23920
rect 66124 23792 66164 27943
rect 66220 27488 66260 28288
rect 66220 27439 66260 27448
rect 66316 25397 66356 28783
rect 66411 26816 66453 26825
rect 66411 26776 66412 26816
rect 66452 26776 66453 26816
rect 66411 26767 66453 26776
rect 66412 25976 66452 26767
rect 66412 25927 66452 25936
rect 66315 25388 66357 25397
rect 66315 25348 66316 25388
rect 66356 25348 66357 25388
rect 66315 25339 66357 25348
rect 66412 25136 66452 25145
rect 66412 24977 66452 25096
rect 66411 24968 66453 24977
rect 66411 24928 66412 24968
rect 66452 24928 66453 24968
rect 66411 24919 66453 24928
rect 66412 24725 66452 24919
rect 66411 24716 66453 24725
rect 66411 24676 66412 24716
rect 66452 24676 66453 24716
rect 66411 24667 66453 24676
rect 66508 23792 66548 23801
rect 66604 23792 66644 31051
rect 66796 29345 66836 31387
rect 66892 31352 66932 32311
rect 66988 31445 67028 34336
rect 67180 34327 67220 34336
rect 67275 34376 67317 34385
rect 67275 34336 67276 34376
rect 67316 34336 67317 34376
rect 67275 34327 67317 34336
rect 67276 34242 67316 34327
rect 67179 34208 67221 34217
rect 67179 34168 67180 34208
rect 67220 34168 67221 34208
rect 67179 34159 67221 34168
rect 67180 33965 67220 34159
rect 67179 33956 67221 33965
rect 67179 33916 67180 33956
rect 67220 33916 67221 33956
rect 67179 33907 67221 33916
rect 67180 32369 67220 33907
rect 67179 32360 67221 32369
rect 67179 32320 67180 32360
rect 67220 32320 67221 32360
rect 67179 32311 67221 32320
rect 67084 32192 67124 32201
rect 67124 32152 67316 32192
rect 67084 32143 67124 32152
rect 67083 31940 67125 31949
rect 67083 31900 67084 31940
rect 67124 31900 67125 31940
rect 67083 31891 67125 31900
rect 66987 31436 67029 31445
rect 66987 31396 66988 31436
rect 67028 31396 67029 31436
rect 66987 31387 67029 31396
rect 66892 31303 66932 31312
rect 67084 31352 67124 31891
rect 67276 31520 67316 32152
rect 67276 31471 67316 31480
rect 66987 31268 67029 31277
rect 66987 31228 66988 31268
rect 67028 31228 67029 31268
rect 66987 31219 67029 31228
rect 66988 31134 67028 31219
rect 67084 31109 67124 31312
rect 67083 31100 67125 31109
rect 67083 31060 67084 31100
rect 67124 31060 67125 31100
rect 67083 31051 67125 31060
rect 67275 30680 67317 30689
rect 67275 30640 67276 30680
rect 67316 30640 67317 30680
rect 67275 30631 67317 30640
rect 67276 29840 67316 30631
rect 67276 29791 67316 29800
rect 66795 29336 66837 29345
rect 66700 29296 66796 29336
rect 66836 29296 66837 29336
rect 66700 25061 66740 29296
rect 66795 29287 66837 29296
rect 66891 28664 66933 28673
rect 66891 28624 66892 28664
rect 66932 28624 66933 28664
rect 66891 28615 66933 28624
rect 66795 28328 66837 28337
rect 66795 28288 66796 28328
rect 66836 28288 66837 28328
rect 66795 28279 66837 28288
rect 66796 27413 66836 28279
rect 66795 27404 66837 27413
rect 66795 27364 66796 27404
rect 66836 27364 66837 27404
rect 66795 27355 66837 27364
rect 66796 26816 66836 27355
rect 66796 25313 66836 26776
rect 66795 25304 66837 25313
rect 66795 25264 66796 25304
rect 66836 25264 66837 25304
rect 66795 25255 66837 25264
rect 66699 25052 66741 25061
rect 66699 25012 66700 25052
rect 66740 25012 66741 25052
rect 66699 25003 66741 25012
rect 66700 24725 66740 25003
rect 66699 24716 66741 24725
rect 66699 24676 66700 24716
rect 66740 24676 66741 24716
rect 66699 24667 66741 24676
rect 66892 23792 66932 28615
rect 67372 28337 67412 34504
rect 67468 34376 67508 34387
rect 67660 34385 67700 34579
rect 67468 34301 67508 34336
rect 67563 34376 67605 34385
rect 67563 34336 67564 34376
rect 67604 34336 67605 34376
rect 67660 34376 67710 34385
rect 67660 34336 67669 34376
rect 67709 34336 67710 34376
rect 67563 34327 67605 34336
rect 67668 34327 67710 34336
rect 67467 34292 67509 34301
rect 67467 34252 67468 34292
rect 67508 34252 67509 34292
rect 67467 34243 67509 34252
rect 67564 34242 67604 34327
rect 67669 34242 67709 34327
rect 67756 34124 67796 36511
rect 67852 35384 67892 37192
rect 68044 35561 68084 37360
rect 68139 37316 68181 37325
rect 68139 37276 68140 37316
rect 68180 37276 68181 37316
rect 68139 37267 68181 37276
rect 68140 36905 68180 37267
rect 68139 36896 68181 36905
rect 68139 36856 68140 36896
rect 68180 36856 68181 36896
rect 68139 36847 68181 36856
rect 68140 36762 68180 36847
rect 68043 35552 68085 35561
rect 68043 35512 68044 35552
rect 68084 35512 68085 35552
rect 68043 35503 68085 35512
rect 67852 35344 68084 35384
rect 67852 35216 67892 35225
rect 67852 34544 67892 35176
rect 68044 34553 68084 35344
rect 68236 35225 68276 37420
rect 68332 37400 68372 37409
rect 68332 37241 68372 37360
rect 68427 37316 68469 37325
rect 68427 37276 68428 37316
rect 68468 37276 68469 37316
rect 68427 37267 68469 37276
rect 68331 37232 68373 37241
rect 68331 37192 68332 37232
rect 68372 37192 68373 37232
rect 68331 37183 68373 37192
rect 68428 37182 68468 37267
rect 68428 36728 68468 36737
rect 68524 36728 68564 38200
rect 68716 37829 68756 38200
rect 68812 38240 68852 38249
rect 68715 37820 68757 37829
rect 68715 37780 68716 37820
rect 68756 37780 68757 37820
rect 68715 37771 68757 37780
rect 68812 37460 68852 38200
rect 69004 38240 69044 38249
rect 70156 38240 70196 38275
rect 69044 38200 69140 38240
rect 69004 38191 69044 38200
rect 69004 37988 69044 37997
rect 69004 37460 69044 37948
rect 69100 37568 69140 38200
rect 70156 38189 70196 38200
rect 71404 38240 71444 38275
rect 72748 38240 72788 38249
rect 71404 38189 71444 38200
rect 72652 38200 72748 38240
rect 69387 38156 69429 38165
rect 69387 38116 69388 38156
rect 69428 38116 69429 38156
rect 69387 38107 69429 38116
rect 70636 38156 70676 38165
rect 69388 38022 69428 38107
rect 69387 37820 69429 37829
rect 69387 37780 69388 37820
rect 69428 37780 69429 37820
rect 69387 37771 69429 37780
rect 69100 37528 69236 37568
rect 68468 36688 68564 36728
rect 68620 37420 68948 37460
rect 69004 37420 69140 37460
rect 68620 36728 68660 37420
rect 68716 37190 68756 37199
rect 68716 36980 68756 37150
rect 68716 36940 68852 36980
rect 68716 36737 68756 36822
rect 68428 36679 68468 36688
rect 68620 36679 68660 36688
rect 68715 36728 68757 36737
rect 68715 36688 68716 36728
rect 68756 36688 68757 36728
rect 68812 36728 68852 36940
rect 68908 36896 68948 37420
rect 69100 37400 69140 37420
rect 69100 37351 69140 37360
rect 69196 37232 69236 37528
rect 69100 37192 69236 37232
rect 69100 36905 69140 37192
rect 69195 36980 69237 36989
rect 69195 36940 69196 36980
rect 69236 36940 69237 36980
rect 69195 36931 69237 36940
rect 69099 36896 69141 36905
rect 68908 36856 69044 36896
rect 69004 36812 69044 36856
rect 69099 36856 69100 36896
rect 69140 36856 69141 36896
rect 69099 36847 69141 36856
rect 69004 36763 69044 36772
rect 68908 36728 68948 36737
rect 68812 36688 68908 36728
rect 68715 36679 68757 36688
rect 68908 36679 68948 36688
rect 69095 36705 69135 36714
rect 69095 36644 69135 36665
rect 69095 36604 69140 36644
rect 68715 36560 68757 36569
rect 68715 36520 68716 36560
rect 68756 36520 68757 36560
rect 68715 36511 68757 36520
rect 68427 36476 68469 36485
rect 68427 36436 68428 36476
rect 68468 36436 68469 36476
rect 68427 36427 68469 36436
rect 68428 36342 68468 36427
rect 68716 36065 68756 36511
rect 69003 36476 69045 36485
rect 69003 36436 69004 36476
rect 69044 36436 69045 36476
rect 69003 36427 69045 36436
rect 68715 36056 68757 36065
rect 68715 36016 68716 36056
rect 68756 36016 68757 36056
rect 68715 36007 68757 36016
rect 68523 35972 68565 35981
rect 68523 35932 68524 35972
rect 68564 35932 68565 35972
rect 68523 35923 68565 35932
rect 68235 35216 68277 35225
rect 68235 35176 68236 35216
rect 68276 35176 68277 35216
rect 68235 35167 68277 35176
rect 67948 34544 67988 34553
rect 67852 34504 67948 34544
rect 67948 34495 67988 34504
rect 68043 34544 68085 34553
rect 68043 34504 68044 34544
rect 68084 34504 68085 34544
rect 68043 34495 68085 34504
rect 67468 34084 67796 34124
rect 67468 33704 67508 34084
rect 67563 33956 67605 33965
rect 67563 33916 67564 33956
rect 67604 33916 67605 33956
rect 67563 33907 67605 33916
rect 67468 33655 67508 33664
rect 67467 29000 67509 29009
rect 67467 28960 67468 29000
rect 67508 28960 67509 29000
rect 67467 28951 67509 28960
rect 67468 28866 67508 28951
rect 66987 28328 67029 28337
rect 66987 28288 66988 28328
rect 67028 28288 67029 28328
rect 66987 28279 67029 28288
rect 67371 28328 67413 28337
rect 67371 28288 67372 28328
rect 67412 28288 67413 28328
rect 67371 28279 67413 28288
rect 66988 28194 67028 28279
rect 67564 27992 67604 33907
rect 67948 32192 67988 32201
rect 67851 31856 67893 31865
rect 67851 31816 67852 31856
rect 67892 31816 67893 31856
rect 67851 31807 67893 31816
rect 67659 29672 67701 29681
rect 67659 29632 67660 29672
rect 67700 29632 67701 29672
rect 67659 29623 67701 29632
rect 67660 29252 67700 29623
rect 67660 29203 67700 29212
rect 67468 27952 67604 27992
rect 67372 27404 67412 27413
rect 67276 27364 67372 27404
rect 67276 26489 67316 27364
rect 67372 27355 67412 27364
rect 67468 27236 67508 27952
rect 67563 27572 67605 27581
rect 67563 27532 67564 27572
rect 67604 27532 67605 27572
rect 67563 27523 67605 27532
rect 67564 27438 67604 27523
rect 67372 27196 67508 27236
rect 67275 26480 67317 26489
rect 67275 26440 67276 26480
rect 67316 26440 67317 26480
rect 67275 26431 67317 26440
rect 67179 26144 67221 26153
rect 67179 26104 67180 26144
rect 67220 26104 67221 26144
rect 67179 26095 67221 26104
rect 67276 26144 67316 26431
rect 67372 26237 67412 27196
rect 67659 26816 67701 26825
rect 67659 26776 67660 26816
rect 67700 26776 67701 26816
rect 67659 26767 67701 26776
rect 67660 26682 67700 26767
rect 67755 26564 67797 26573
rect 67755 26524 67756 26564
rect 67796 26524 67797 26564
rect 67755 26515 67797 26524
rect 67756 26312 67796 26515
rect 67852 26321 67892 31807
rect 67948 30689 67988 32152
rect 67947 30680 67989 30689
rect 67947 30640 67948 30680
rect 67988 30640 67989 30680
rect 67947 30631 67989 30640
rect 68236 30680 68276 30689
rect 68236 29765 68276 30640
rect 68331 29840 68373 29849
rect 68331 29800 68332 29840
rect 68372 29800 68373 29840
rect 68331 29791 68373 29800
rect 68235 29756 68277 29765
rect 68235 29716 68236 29756
rect 68276 29716 68277 29756
rect 68235 29707 68277 29716
rect 68332 29672 68372 29791
rect 68428 29672 68468 29681
rect 68332 29632 68428 29672
rect 68044 29168 68084 29177
rect 68044 29009 68084 29128
rect 68043 29000 68085 29009
rect 68043 28960 68044 29000
rect 68084 28960 68085 29000
rect 68043 28951 68085 28960
rect 68332 28841 68372 29632
rect 68428 29623 68468 29632
rect 68427 29252 68469 29261
rect 68427 29212 68428 29252
rect 68468 29212 68469 29252
rect 68427 29203 68469 29212
rect 68331 28832 68373 28841
rect 68331 28792 68332 28832
rect 68372 28792 68373 28832
rect 68331 28783 68373 28792
rect 68140 28160 68180 28171
rect 68140 28085 68180 28120
rect 68139 28076 68181 28085
rect 68139 28036 68140 28076
rect 68180 28036 68181 28076
rect 68139 28027 68181 28036
rect 68140 27665 68180 28027
rect 68139 27656 68181 27665
rect 68139 27616 68140 27656
rect 68180 27616 68181 27656
rect 68139 27607 68181 27616
rect 68331 27488 68373 27497
rect 68331 27448 68332 27488
rect 68372 27448 68373 27488
rect 68331 27439 68373 27448
rect 68332 26816 68372 27439
rect 68428 26825 68468 29203
rect 68524 27572 68564 35923
rect 68716 35216 68756 36007
rect 68811 35720 68853 35729
rect 68811 35680 68812 35720
rect 68852 35680 68853 35720
rect 68811 35671 68853 35680
rect 68716 35167 68756 35176
rect 68620 33452 68660 33461
rect 68620 32873 68660 33412
rect 68812 33140 68852 35671
rect 68907 34628 68949 34637
rect 68907 34588 68908 34628
rect 68948 34588 68949 34628
rect 68907 34579 68949 34588
rect 68908 34494 68948 34579
rect 69004 34469 69044 36427
rect 69100 36401 69140 36604
rect 69196 36560 69236 36931
rect 69291 36896 69333 36905
rect 69291 36856 69292 36896
rect 69332 36856 69333 36896
rect 69291 36847 69333 36856
rect 69292 36728 69332 36847
rect 69388 36812 69428 37771
rect 69484 37400 69524 37409
rect 70348 37400 70388 37409
rect 70636 37400 70676 38116
rect 69524 37360 69716 37400
rect 69484 37351 69524 37360
rect 69483 37232 69525 37241
rect 69483 37192 69484 37232
rect 69524 37192 69525 37232
rect 69483 37183 69525 37192
rect 69484 36821 69524 37183
rect 69388 36763 69428 36772
rect 69483 36812 69525 36821
rect 69483 36772 69484 36812
rect 69524 36772 69525 36812
rect 69483 36763 69525 36772
rect 69292 36679 69332 36688
rect 69484 36728 69524 36763
rect 69484 36677 69524 36688
rect 69676 36560 69716 37360
rect 70388 37360 70676 37400
rect 70348 37351 70388 37360
rect 70539 36896 70581 36905
rect 70539 36856 70540 36896
rect 70580 36856 70581 36896
rect 70539 36847 70581 36856
rect 69771 36728 69813 36737
rect 69771 36688 69772 36728
rect 69812 36688 69813 36728
rect 69771 36679 69813 36688
rect 69196 36520 69428 36560
rect 69099 36392 69141 36401
rect 69099 36352 69100 36392
rect 69140 36352 69141 36392
rect 69099 36343 69141 36352
rect 69099 36224 69141 36233
rect 69099 36184 69100 36224
rect 69140 36184 69141 36224
rect 69099 36175 69141 36184
rect 69003 34460 69045 34469
rect 69003 34420 69004 34460
rect 69044 34420 69045 34460
rect 69003 34411 69045 34420
rect 68716 33100 68852 33140
rect 68619 32864 68661 32873
rect 68619 32824 68620 32864
rect 68660 32824 68661 32864
rect 68619 32815 68661 32824
rect 68619 31520 68661 31529
rect 68619 31480 68620 31520
rect 68660 31480 68661 31520
rect 68619 31471 68661 31480
rect 68620 30680 68660 31471
rect 68620 30631 68660 30640
rect 68716 30596 68756 33100
rect 68811 32864 68853 32873
rect 68811 32824 68812 32864
rect 68852 32824 68853 32864
rect 68811 32815 68853 32824
rect 68908 32864 68948 32873
rect 68812 32730 68852 32815
rect 68908 32453 68948 32824
rect 69100 32864 69140 36175
rect 69195 34880 69237 34889
rect 69195 34840 69196 34880
rect 69236 34840 69237 34880
rect 69195 34831 69237 34840
rect 69003 32696 69045 32705
rect 69003 32656 69004 32696
rect 69044 32656 69045 32696
rect 69003 32647 69045 32656
rect 69004 32562 69044 32647
rect 69100 32537 69140 32824
rect 69099 32528 69141 32537
rect 69099 32488 69100 32528
rect 69140 32488 69141 32528
rect 69099 32479 69141 32488
rect 68907 32444 68949 32453
rect 68907 32404 68908 32444
rect 68948 32404 69044 32444
rect 68907 32395 68949 32404
rect 68811 31520 68853 31529
rect 68811 31480 68812 31520
rect 68852 31480 68853 31520
rect 68811 31471 68853 31480
rect 68812 31386 68852 31471
rect 68907 30680 68949 30689
rect 68907 30640 68908 30680
rect 68948 30640 68949 30680
rect 68907 30631 68949 30640
rect 68716 30556 68852 30596
rect 68524 27532 68756 27572
rect 68523 27404 68565 27413
rect 68523 27364 68524 27404
rect 68564 27364 68565 27404
rect 68523 27355 68565 27364
rect 68332 26767 68372 26776
rect 68427 26816 68469 26825
rect 68427 26776 68428 26816
rect 68468 26776 68469 26816
rect 68427 26767 68469 26776
rect 68524 26816 68564 27355
rect 68044 26732 68084 26741
rect 68044 26573 68084 26692
rect 68428 26648 68468 26657
rect 68332 26608 68428 26648
rect 68043 26564 68085 26573
rect 68043 26524 68044 26564
rect 68084 26524 68085 26564
rect 68043 26515 68085 26524
rect 68332 26396 68372 26608
rect 68428 26599 68468 26608
rect 67948 26356 68372 26396
rect 68427 26396 68469 26405
rect 68427 26356 68428 26396
rect 68468 26356 68469 26396
rect 67756 26263 67796 26272
rect 67851 26312 67893 26321
rect 67851 26272 67852 26312
rect 67892 26272 67893 26312
rect 67851 26263 67893 26272
rect 67371 26228 67413 26237
rect 67371 26188 67372 26228
rect 67412 26188 67413 26228
rect 67371 26179 67413 26188
rect 67276 26095 67316 26104
rect 67372 26144 67412 26179
rect 67180 25976 67220 26095
rect 67372 26094 67412 26104
rect 67468 26144 67508 26153
rect 67660 26144 67700 26153
rect 67508 26104 67660 26144
rect 67468 26095 67508 26104
rect 67660 26095 67700 26104
rect 67852 26144 67892 26153
rect 67180 25936 67508 25976
rect 67083 25388 67125 25397
rect 67083 25348 67084 25388
rect 67124 25348 67125 25388
rect 67083 25339 67125 25348
rect 67084 25304 67124 25339
rect 67084 25253 67124 25264
rect 67372 25304 67412 25313
rect 67372 24809 67412 25264
rect 67468 25304 67508 25936
rect 67852 25901 67892 26104
rect 67948 26144 67988 26356
rect 68427 26347 68469 26356
rect 67948 26095 67988 26104
rect 68140 26144 68180 26153
rect 67851 25892 67893 25901
rect 67851 25852 67852 25892
rect 67892 25852 67893 25892
rect 67851 25843 67893 25852
rect 67852 25724 67892 25843
rect 68140 25733 68180 26104
rect 68332 26144 68372 26153
rect 68235 25892 68277 25901
rect 68235 25852 68236 25892
rect 68276 25852 68277 25892
rect 68235 25843 68277 25852
rect 68236 25758 68276 25843
rect 67468 25255 67508 25264
rect 67660 25684 67892 25724
rect 68139 25724 68181 25733
rect 68139 25684 68140 25724
rect 68180 25684 68181 25724
rect 67660 25061 67700 25684
rect 68139 25675 68181 25684
rect 67756 25556 67796 25565
rect 68332 25556 68372 26104
rect 67796 25516 68372 25556
rect 67756 25507 67796 25516
rect 68428 25388 68468 26347
rect 68524 25976 68564 26776
rect 68620 26816 68660 26825
rect 68620 26153 68660 26776
rect 68619 26144 68661 26153
rect 68619 26104 68620 26144
rect 68660 26104 68661 26144
rect 68619 26095 68661 26104
rect 68620 25976 68660 25985
rect 68524 25936 68620 25976
rect 68620 25927 68660 25936
rect 68428 25348 68660 25388
rect 68332 25291 68372 25300
rect 67948 25220 67988 25229
rect 67756 25180 67948 25220
rect 67659 25052 67701 25061
rect 67659 25012 67660 25052
rect 67700 25012 67701 25052
rect 67659 25003 67701 25012
rect 67371 24800 67413 24809
rect 67371 24760 67372 24800
rect 67412 24760 67413 24800
rect 67371 24751 67413 24760
rect 67756 24800 67796 25180
rect 67948 25171 67988 25180
rect 68332 25136 68372 25251
rect 68332 25096 68564 25136
rect 67851 25052 67893 25061
rect 67851 25012 67852 25052
rect 67892 25012 67893 25052
rect 67851 25003 67893 25012
rect 67756 24751 67796 24760
rect 67659 24716 67701 24725
rect 67659 24676 67660 24716
rect 67700 24676 67701 24716
rect 67659 24667 67701 24676
rect 67660 24632 67700 24667
rect 67660 24581 67700 24592
rect 67852 24632 67892 25003
rect 68331 24800 68373 24809
rect 67852 24583 67892 24592
rect 67948 24760 68276 24800
rect 67948 24632 67988 24760
rect 68236 24716 68276 24760
rect 68331 24760 68332 24800
rect 68372 24760 68373 24800
rect 68331 24751 68373 24760
rect 68236 24667 68276 24676
rect 67948 24583 67988 24592
rect 68139 24632 68181 24641
rect 68139 24592 68140 24632
rect 68180 24592 68181 24632
rect 68139 24583 68181 24592
rect 68332 24632 68372 24751
rect 68332 24583 68372 24592
rect 67275 24548 67317 24557
rect 67275 24508 67276 24548
rect 67316 24508 67317 24548
rect 67275 24499 67317 24508
rect 67276 23801 67316 24499
rect 68140 24498 68180 24583
rect 68524 24464 68564 25096
rect 68524 24415 68564 24424
rect 68620 24296 68660 25348
rect 68140 24256 68660 24296
rect 67755 24044 67797 24053
rect 67755 24004 67756 24044
rect 67796 24004 67797 24044
rect 67755 23995 67797 24004
rect 67275 23792 67317 23801
rect 65780 23752 66068 23792
rect 65740 23743 65780 23752
rect 65836 23624 65876 23633
rect 65836 23060 65876 23584
rect 66028 23060 66068 23752
rect 66164 23752 66452 23792
rect 66124 23743 66164 23752
rect 66220 23624 66260 23633
rect 66220 23060 66260 23584
rect 66412 23060 66452 23752
rect 66548 23752 66836 23792
rect 66508 23743 66548 23752
rect 66604 23624 66644 23633
rect 66604 23060 66644 23584
rect 66796 23060 66836 23752
rect 66932 23752 67220 23792
rect 66892 23743 66932 23752
rect 66988 23624 67028 23633
rect 66988 23060 67028 23584
rect 67180 23060 67220 23752
rect 67275 23752 67276 23792
rect 67316 23752 67317 23792
rect 67275 23743 67317 23752
rect 67659 23792 67701 23801
rect 67659 23752 67660 23792
rect 67700 23752 67701 23792
rect 67659 23743 67701 23752
rect 67756 23792 67796 23995
rect 68140 23792 68180 24256
rect 67796 23752 68084 23792
rect 67756 23743 67796 23752
rect 67276 23658 67316 23743
rect 67372 23624 67412 23633
rect 67372 23060 67412 23584
rect 65356 23020 65585 23060
rect 65644 23020 65695 23060
rect 65836 23020 65985 23060
rect 66028 23020 66095 23060
rect 66220 23020 66356 23060
rect 66412 23020 66495 23060
rect 66604 23020 66740 23060
rect 66796 23020 66895 23060
rect 66988 23020 67124 23060
rect 67180 23020 67295 23060
rect 67372 23020 67508 23060
rect 65255 22596 65295 23020
rect 65545 22596 65585 23020
rect 65655 22596 65695 23020
rect 65945 22596 65985 23020
rect 66055 22596 66095 23020
rect 66316 22784 66356 23020
rect 66316 22744 66385 22784
rect 66345 22596 66385 22744
rect 66455 22596 66495 23020
rect 66700 22784 66740 23020
rect 66700 22744 66785 22784
rect 66745 22596 66785 22744
rect 66855 22596 66895 23020
rect 67084 22784 67124 23020
rect 67084 22744 67185 22784
rect 67145 22596 67185 22744
rect 67255 22596 67295 23020
rect 67468 22784 67508 23020
rect 67660 22784 67700 23743
rect 67468 22744 67585 22784
rect 67545 22596 67585 22744
rect 67655 22744 67700 22784
rect 67852 23624 67892 23633
rect 67852 22784 67892 23584
rect 68044 23060 68084 23752
rect 68140 23743 68180 23752
rect 68236 23624 68276 23633
rect 68236 23060 68276 23584
rect 68428 23060 68468 24256
rect 68523 23960 68565 23969
rect 68523 23920 68524 23960
rect 68564 23920 68565 23960
rect 68523 23911 68565 23920
rect 68524 23792 68564 23911
rect 68716 23801 68756 27532
rect 68812 27245 68852 30556
rect 68908 29168 68948 30631
rect 69004 30092 69044 32404
rect 69100 31940 69140 31949
rect 69100 31109 69140 31900
rect 69099 31100 69141 31109
rect 69099 31060 69100 31100
rect 69140 31060 69141 31100
rect 69099 31051 69141 31060
rect 69100 30092 69140 30101
rect 69004 30052 69100 30092
rect 69100 29849 69140 30052
rect 69099 29840 69141 29849
rect 69099 29800 69100 29840
rect 69140 29800 69141 29840
rect 69099 29791 69141 29800
rect 68908 29119 68948 29128
rect 68907 27908 68949 27917
rect 68907 27868 68908 27908
rect 68948 27868 68949 27908
rect 68907 27859 68949 27868
rect 68908 27497 68948 27859
rect 69196 27740 69236 34831
rect 69292 32780 69332 32789
rect 69292 32369 69332 32740
rect 69291 32360 69333 32369
rect 69291 32320 69292 32360
rect 69332 32320 69333 32360
rect 69291 32311 69333 32320
rect 69291 30008 69333 30017
rect 69291 29968 69292 30008
rect 69332 29968 69333 30008
rect 69291 29959 69333 29968
rect 69292 29924 69332 29959
rect 69292 29873 69332 29884
rect 69388 27833 69428 36520
rect 69676 36511 69716 36520
rect 69675 36224 69717 36233
rect 69675 36184 69676 36224
rect 69716 36184 69717 36224
rect 69675 36175 69717 36184
rect 69483 36140 69525 36149
rect 69483 36100 69484 36140
rect 69524 36100 69525 36140
rect 69483 36091 69525 36100
rect 69484 36056 69524 36091
rect 69484 36005 69524 36016
rect 69676 35888 69716 36175
rect 69676 35839 69716 35848
rect 69772 35804 69812 36679
rect 70059 36560 70101 36569
rect 70059 36520 70060 36560
rect 70100 36520 70101 36560
rect 70059 36511 70101 36520
rect 70060 36065 70100 36511
rect 70059 36056 70101 36065
rect 70059 36016 70060 36056
rect 70100 36016 70101 36056
rect 70059 36007 70101 36016
rect 69867 35888 69909 35897
rect 69867 35848 69868 35888
rect 69908 35848 69909 35888
rect 69867 35839 69909 35848
rect 69964 35888 70004 35897
rect 69772 35755 69812 35764
rect 69868 35754 69908 35839
rect 69868 34964 69908 34973
rect 69868 34385 69908 34924
rect 69964 34637 70004 35848
rect 69963 34628 70005 34637
rect 69963 34588 69964 34628
rect 70004 34588 70005 34628
rect 69963 34579 70005 34588
rect 69867 34376 69909 34385
rect 69867 34336 69868 34376
rect 69908 34336 69909 34376
rect 69867 34327 69909 34336
rect 70060 34376 70100 36007
rect 70540 35477 70580 36847
rect 70636 36569 70676 37360
rect 71980 38072 72020 38081
rect 71115 37232 71157 37241
rect 71115 37192 71116 37232
rect 71156 37192 71157 37232
rect 71115 37183 71157 37192
rect 71499 37232 71541 37241
rect 71499 37192 71500 37232
rect 71540 37192 71541 37232
rect 71499 37183 71541 37192
rect 71116 36821 71156 37183
rect 71500 37098 71540 37183
rect 71980 37073 72020 38032
rect 71979 37064 72021 37073
rect 71979 37024 71980 37064
rect 72020 37024 72021 37064
rect 71979 37015 72021 37024
rect 71115 36812 71157 36821
rect 71115 36772 71116 36812
rect 71156 36772 71157 36812
rect 71115 36763 71157 36772
rect 70635 36560 70677 36569
rect 70635 36520 70636 36560
rect 70676 36520 70677 36560
rect 70635 36511 70677 36520
rect 70923 36476 70965 36485
rect 70923 36436 70924 36476
rect 70964 36436 70965 36476
rect 70923 36427 70965 36436
rect 70924 36342 70964 36427
rect 70923 36140 70965 36149
rect 70923 36100 70924 36140
rect 70964 36100 70965 36140
rect 70923 36091 70965 36100
rect 70539 35468 70581 35477
rect 70539 35428 70540 35468
rect 70580 35428 70581 35468
rect 70539 35419 70581 35428
rect 70827 35468 70869 35477
rect 70827 35428 70828 35468
rect 70868 35428 70869 35468
rect 70827 35419 70869 35428
rect 70444 35309 70484 35340
rect 70443 35300 70485 35309
rect 70443 35260 70444 35300
rect 70484 35260 70485 35300
rect 70443 35251 70485 35260
rect 70444 35216 70484 35251
rect 70444 34637 70484 35176
rect 70539 35216 70581 35225
rect 70539 35176 70540 35216
rect 70580 35176 70581 35216
rect 70539 35167 70581 35176
rect 70636 35216 70676 35225
rect 70443 34628 70485 34637
rect 70443 34588 70444 34628
rect 70484 34588 70485 34628
rect 70443 34579 70485 34588
rect 70347 34544 70389 34553
rect 70347 34504 70348 34544
rect 70388 34504 70389 34544
rect 70347 34495 70389 34504
rect 70060 34327 70100 34336
rect 69579 34124 69621 34133
rect 69579 34084 69580 34124
rect 69620 34084 69621 34124
rect 69579 34075 69621 34084
rect 69483 31688 69525 31697
rect 69483 31648 69484 31688
rect 69524 31648 69525 31688
rect 69483 31639 69525 31648
rect 69484 30689 69524 31639
rect 69483 30680 69525 30689
rect 69483 30640 69484 30680
rect 69524 30640 69525 30680
rect 69483 30631 69525 30640
rect 69484 30546 69524 30631
rect 69483 30092 69525 30101
rect 69483 30052 69484 30092
rect 69524 30052 69525 30092
rect 69483 30043 69525 30052
rect 69484 29924 69524 30043
rect 69484 27917 69524 29884
rect 69483 27908 69525 27917
rect 69483 27868 69484 27908
rect 69524 27868 69525 27908
rect 69580 27908 69620 34075
rect 69868 33965 69908 34327
rect 69867 33956 69909 33965
rect 69867 33916 69868 33956
rect 69908 33916 69909 33956
rect 69867 33907 69909 33916
rect 69772 33536 69812 33545
rect 69676 33496 69772 33536
rect 69676 32864 69716 33496
rect 69772 33487 69812 33496
rect 70348 33209 70388 34495
rect 70347 33200 70389 33209
rect 70347 33160 70348 33200
rect 70388 33160 70389 33200
rect 70347 33151 70389 33160
rect 69676 32815 69716 32824
rect 69771 32696 69813 32705
rect 69771 32656 69772 32696
rect 69812 32656 69813 32696
rect 69771 32647 69813 32656
rect 69675 32528 69717 32537
rect 69675 32488 69676 32528
rect 69716 32488 69717 32528
rect 69675 32479 69717 32488
rect 69676 30092 69716 32479
rect 69772 32192 69812 32647
rect 69963 32360 70005 32369
rect 69963 32320 69964 32360
rect 70004 32320 70005 32360
rect 69963 32311 70005 32320
rect 69964 32226 70004 32311
rect 69772 32143 69812 32152
rect 69868 32192 69908 32201
rect 69868 32033 69908 32152
rect 70060 32192 70100 32201
rect 70252 32192 70292 32201
rect 70100 32152 70252 32192
rect 70060 32143 70100 32152
rect 70252 32143 70292 32152
rect 70348 32192 70388 33151
rect 70540 33140 70580 35167
rect 70636 34553 70676 35176
rect 70731 35216 70773 35225
rect 70731 35176 70732 35216
rect 70772 35176 70773 35216
rect 70731 35167 70773 35176
rect 70732 35082 70772 35167
rect 70635 34544 70677 34553
rect 70635 34504 70636 34544
rect 70676 34504 70677 34544
rect 70635 34495 70677 34504
rect 70828 33140 70868 35419
rect 70924 34376 70964 36091
rect 71019 35552 71061 35561
rect 71019 35512 71020 35552
rect 71060 35512 71061 35552
rect 71019 35503 71061 35512
rect 70924 34327 70964 34336
rect 71020 35216 71060 35503
rect 69867 32024 69909 32033
rect 69867 31984 69868 32024
rect 69908 31984 69909 32024
rect 69867 31975 69909 31984
rect 70348 31352 70388 32152
rect 70444 33100 70580 33140
rect 70732 33100 70868 33140
rect 70444 32192 70484 33100
rect 70540 32864 70580 32873
rect 70580 32824 70676 32864
rect 70540 32815 70580 32824
rect 70539 32696 70581 32705
rect 70539 32656 70540 32696
rect 70580 32656 70581 32696
rect 70539 32647 70581 32656
rect 70444 31520 70484 32152
rect 70540 32192 70580 32647
rect 70540 32143 70580 32152
rect 70636 31697 70676 32824
rect 70635 31688 70677 31697
rect 70635 31648 70636 31688
rect 70676 31648 70677 31688
rect 70635 31639 70677 31648
rect 70732 31613 70772 33100
rect 70827 32696 70869 32705
rect 70827 32656 70828 32696
rect 70868 32656 70869 32696
rect 70827 32647 70869 32656
rect 70828 32192 70868 32647
rect 70923 32444 70965 32453
rect 70923 32404 70924 32444
rect 70964 32404 70965 32444
rect 70923 32395 70965 32404
rect 70828 32143 70868 32152
rect 70924 32192 70964 32395
rect 71020 32369 71060 35176
rect 71116 32957 71156 36763
rect 72076 36728 72116 36737
rect 72076 36569 72116 36688
rect 72075 36560 72117 36569
rect 72075 36520 72076 36560
rect 72116 36520 72117 36560
rect 72075 36511 72117 36520
rect 72171 36476 72213 36485
rect 72171 36436 72172 36476
rect 72212 36436 72213 36476
rect 72171 36427 72213 36436
rect 71211 36140 71253 36149
rect 71211 36100 71212 36140
rect 71252 36100 71253 36140
rect 71211 36091 71253 36100
rect 71883 36140 71925 36149
rect 71883 36100 71884 36140
rect 71924 36100 71925 36140
rect 71883 36091 71925 36100
rect 71115 32948 71157 32957
rect 71115 32908 71116 32948
rect 71156 32908 71157 32948
rect 71115 32899 71157 32908
rect 71115 32528 71157 32537
rect 71115 32488 71116 32528
rect 71156 32488 71157 32528
rect 71115 32479 71157 32488
rect 71019 32360 71061 32369
rect 71019 32320 71020 32360
rect 71060 32320 71061 32360
rect 71019 32311 71061 32320
rect 71116 32285 71156 32479
rect 71115 32276 71157 32285
rect 71115 32236 71116 32276
rect 71156 32236 71157 32276
rect 71115 32227 71157 32236
rect 70924 32143 70964 32152
rect 71116 32192 71156 32227
rect 71116 32141 71156 32152
rect 71116 31940 71156 31949
rect 71020 31900 71116 31940
rect 70731 31604 70773 31613
rect 70731 31564 70732 31604
rect 70772 31564 70773 31604
rect 70731 31555 70773 31564
rect 70444 31480 70676 31520
rect 70540 31352 70580 31361
rect 70348 31312 70540 31352
rect 70443 31184 70485 31193
rect 70443 31144 70444 31184
rect 70484 31144 70485 31184
rect 70443 31135 70485 31144
rect 70444 31050 70484 31135
rect 70540 30932 70580 31312
rect 70636 31352 70676 31480
rect 70923 31436 70965 31445
rect 70923 31396 70924 31436
rect 70964 31396 70965 31436
rect 70923 31387 70965 31396
rect 70636 31100 70676 31312
rect 70731 31352 70773 31361
rect 70731 31312 70732 31352
rect 70772 31312 70773 31352
rect 70731 31303 70773 31312
rect 70732 31218 70772 31303
rect 70924 31302 70964 31387
rect 70827 31184 70869 31193
rect 70827 31144 70828 31184
rect 70868 31144 70869 31184
rect 70827 31135 70869 31144
rect 70636 31060 70785 31100
rect 70745 30932 70785 31060
rect 69676 30043 69716 30052
rect 70444 30892 70580 30932
rect 70732 30892 70785 30932
rect 70348 30008 70388 30017
rect 70156 29968 70348 30008
rect 69868 29840 69908 29849
rect 69676 29672 69716 29681
rect 69676 29588 69716 29632
rect 69771 29588 69813 29597
rect 69676 29548 69772 29588
rect 69812 29548 69813 29588
rect 69771 29539 69813 29548
rect 69868 29336 69908 29800
rect 70060 29840 70100 29849
rect 69963 29672 70005 29681
rect 69963 29632 69964 29672
rect 70004 29632 70005 29672
rect 69963 29623 70005 29632
rect 69964 29538 70004 29623
rect 70060 29513 70100 29800
rect 70156 29840 70196 29968
rect 70348 29959 70388 29968
rect 70348 29840 70388 29849
rect 70156 29791 70196 29800
rect 70252 29800 70348 29840
rect 70252 29597 70292 29800
rect 70348 29791 70388 29800
rect 70444 29672 70484 30892
rect 70635 30764 70677 30773
rect 70635 30724 70636 30764
rect 70676 30724 70677 30764
rect 70635 30715 70677 30724
rect 70539 30680 70581 30689
rect 70539 30640 70540 30680
rect 70580 30640 70581 30680
rect 70539 30631 70581 30640
rect 70540 30101 70580 30631
rect 70636 30428 70676 30715
rect 70539 30092 70581 30101
rect 70539 30052 70540 30092
rect 70580 30052 70581 30092
rect 70539 30043 70581 30052
rect 70539 29840 70581 29849
rect 70539 29800 70540 29840
rect 70580 29800 70581 29840
rect 70539 29791 70581 29800
rect 70636 29840 70676 30388
rect 70732 30101 70772 30892
rect 70731 30092 70773 30101
rect 70731 30052 70732 30092
rect 70772 30052 70773 30092
rect 70731 30043 70773 30052
rect 70636 29791 70676 29800
rect 70540 29706 70580 29791
rect 70348 29632 70484 29672
rect 70251 29588 70293 29597
rect 70251 29548 70252 29588
rect 70292 29548 70293 29588
rect 70251 29539 70293 29548
rect 70059 29504 70101 29513
rect 70059 29464 70060 29504
rect 70100 29464 70101 29504
rect 70059 29455 70101 29464
rect 70252 29336 70292 29345
rect 69868 29296 70252 29336
rect 70252 29287 70292 29296
rect 70348 29168 70388 29632
rect 70635 29504 70677 29513
rect 70635 29464 70636 29504
rect 70676 29464 70677 29504
rect 70635 29455 70677 29464
rect 70348 29119 70388 29128
rect 70443 29168 70485 29177
rect 70443 29128 70444 29168
rect 70484 29128 70485 29168
rect 70443 29119 70485 29128
rect 70540 29168 70580 29179
rect 70059 29084 70101 29093
rect 70059 29044 70060 29084
rect 70100 29044 70101 29084
rect 70059 29035 70101 29044
rect 70060 28950 70100 29035
rect 70444 29034 70484 29119
rect 70540 29093 70580 29128
rect 70539 29084 70581 29093
rect 70539 29044 70540 29084
rect 70580 29044 70581 29084
rect 70539 29035 70581 29044
rect 70251 29000 70293 29009
rect 70251 28960 70252 29000
rect 70292 28960 70293 29000
rect 70251 28951 70293 28960
rect 70252 28328 70292 28951
rect 70540 28496 70580 29035
rect 70636 28580 70676 29455
rect 70732 29336 70772 30043
rect 70828 29840 70868 31135
rect 71020 30848 71060 31900
rect 71116 31891 71156 31900
rect 71115 31604 71157 31613
rect 71115 31564 71116 31604
rect 71156 31564 71157 31604
rect 71115 31555 71157 31564
rect 71116 31470 71156 31555
rect 71115 31184 71157 31193
rect 71115 31144 71116 31184
rect 71156 31144 71157 31184
rect 71115 31135 71157 31144
rect 71116 31050 71156 31135
rect 71212 30857 71252 36091
rect 71595 35888 71637 35897
rect 71595 35848 71596 35888
rect 71636 35848 71637 35888
rect 71595 35839 71637 35848
rect 71884 35888 71924 36091
rect 71884 35839 71924 35848
rect 71979 35888 72021 35897
rect 72172 35888 72212 36427
rect 72555 36392 72597 36401
rect 72555 36352 72556 36392
rect 72596 36352 72597 36392
rect 72555 36343 72597 36352
rect 71979 35848 71980 35888
rect 72020 35874 72116 35888
rect 72020 35848 72076 35874
rect 71979 35839 72021 35848
rect 71403 35300 71445 35309
rect 71403 35260 71404 35300
rect 71444 35260 71445 35300
rect 71403 35251 71445 35260
rect 71308 35216 71348 35225
rect 71308 34712 71348 35176
rect 71404 35166 71444 35251
rect 71308 34672 71444 34712
rect 71307 34544 71349 34553
rect 71307 34504 71308 34544
rect 71348 34504 71349 34544
rect 71307 34495 71349 34504
rect 71308 34376 71348 34495
rect 71308 34327 71348 34336
rect 71404 34217 71444 34672
rect 71403 34208 71445 34217
rect 71403 34168 71404 34208
rect 71444 34168 71445 34208
rect 71403 34159 71445 34168
rect 71596 33713 71636 35839
rect 72172 35839 72212 35848
rect 72076 35825 72116 35834
rect 71980 35720 72020 35729
rect 72020 35680 72212 35720
rect 71980 35671 72020 35680
rect 71883 35216 71925 35225
rect 71883 35176 71884 35216
rect 71924 35176 71925 35216
rect 71883 35167 71925 35176
rect 72076 35216 72116 35225
rect 71884 35082 71924 35167
rect 71691 35048 71733 35057
rect 71691 35008 71692 35048
rect 71732 35008 71733 35048
rect 71691 34999 71733 35008
rect 71692 34914 71732 34999
rect 72076 34973 72116 35176
rect 72172 35216 72212 35680
rect 72556 35309 72596 36343
rect 72555 35300 72597 35309
rect 72555 35260 72556 35300
rect 72596 35260 72597 35300
rect 72555 35251 72597 35260
rect 72172 35167 72212 35176
rect 72364 35216 72404 35225
rect 72364 35057 72404 35176
rect 72556 35216 72596 35251
rect 72556 35166 72596 35176
rect 72363 35048 72405 35057
rect 72363 35008 72364 35048
rect 72404 35008 72405 35048
rect 72363 34999 72405 35008
rect 72555 35048 72597 35057
rect 72555 35008 72556 35048
rect 72596 35008 72597 35048
rect 72555 34999 72597 35008
rect 71884 34964 71924 34973
rect 71788 34924 71884 34964
rect 71788 34553 71828 34924
rect 71884 34915 71924 34924
rect 72075 34964 72117 34973
rect 72075 34924 72076 34964
rect 72116 34924 72117 34964
rect 72075 34915 72117 34924
rect 72459 34964 72501 34973
rect 72459 34924 72460 34964
rect 72500 34924 72501 34964
rect 72459 34915 72501 34924
rect 72076 34796 72116 34915
rect 72460 34830 72500 34915
rect 71884 34756 72116 34796
rect 71787 34544 71829 34553
rect 71787 34504 71788 34544
rect 71828 34504 71829 34544
rect 71787 34495 71829 34504
rect 71692 34376 71732 34385
rect 71692 33788 71732 34336
rect 71788 34376 71828 34385
rect 71884 34376 71924 34756
rect 71980 34544 72020 34553
rect 72020 34504 72212 34544
rect 71980 34495 72020 34504
rect 71828 34336 71924 34376
rect 71979 34376 72021 34385
rect 71979 34336 71980 34376
rect 72020 34336 72021 34376
rect 71788 34327 71828 34336
rect 71979 34327 72021 34336
rect 72172 34376 72212 34504
rect 72172 34327 72212 34336
rect 72556 34376 72596 34999
rect 72556 34327 72596 34336
rect 71787 34208 71829 34217
rect 71787 34168 71788 34208
rect 71828 34168 71829 34208
rect 71787 34159 71829 34168
rect 71692 33739 71732 33748
rect 71595 33704 71637 33713
rect 71500 33664 71596 33704
rect 71636 33664 71637 33704
rect 71500 32453 71540 33664
rect 71595 33655 71637 33664
rect 71788 33704 71828 34159
rect 71980 33881 72020 34327
rect 72652 33956 72692 38200
rect 72748 38191 72788 38200
rect 76876 38240 76916 38249
rect 77164 38240 77204 38249
rect 76916 38200 77012 38240
rect 76876 38191 76916 38200
rect 73996 38072 74036 38081
rect 76012 38072 76052 38081
rect 74036 38032 74132 38072
rect 73996 38023 74036 38032
rect 73036 37988 73076 37997
rect 73076 37948 73172 37988
rect 73036 37939 73076 37948
rect 73036 37493 73076 37524
rect 73035 37484 73077 37493
rect 73035 37444 73036 37484
rect 73076 37444 73077 37484
rect 73035 37435 73077 37444
rect 72748 37400 72788 37409
rect 72748 36485 72788 37360
rect 72844 37400 72884 37409
rect 72844 36737 72884 37360
rect 72940 37400 72980 37409
rect 72940 37241 72980 37360
rect 73036 37316 73076 37435
rect 73036 37267 73076 37276
rect 72939 37232 72981 37241
rect 72939 37192 72940 37232
rect 72980 37192 72981 37232
rect 72939 37183 72981 37192
rect 72939 37064 72981 37073
rect 72939 37024 72940 37064
rect 72980 37024 72981 37064
rect 72939 37015 72981 37024
rect 72843 36728 72885 36737
rect 72843 36688 72844 36728
rect 72884 36688 72885 36728
rect 72843 36679 72885 36688
rect 72940 36728 72980 37015
rect 72940 36679 72980 36688
rect 72747 36476 72789 36485
rect 72747 36436 72748 36476
rect 72788 36436 72789 36476
rect 72747 36427 72789 36436
rect 72748 35888 72788 35897
rect 72748 35225 72788 35848
rect 72747 35216 72789 35225
rect 72747 35176 72748 35216
rect 72788 35176 72789 35216
rect 72747 35167 72789 35176
rect 72747 35048 72789 35057
rect 72747 35008 72748 35048
rect 72788 35008 72789 35048
rect 72747 34999 72789 35008
rect 72748 34914 72788 34999
rect 72652 33916 72788 33956
rect 71979 33872 72021 33881
rect 71979 33832 71980 33872
rect 72020 33832 72021 33872
rect 71979 33823 72021 33832
rect 71980 33704 72020 33823
rect 72172 33704 72212 33713
rect 71788 33655 71828 33664
rect 71884 33664 71980 33704
rect 71596 33570 71636 33655
rect 71884 33140 71924 33664
rect 71980 33655 72020 33664
rect 72076 33664 72172 33704
rect 71788 33100 71924 33140
rect 71980 33452 72020 33461
rect 71691 32696 71733 32705
rect 71691 32656 71692 32696
rect 71732 32656 71733 32696
rect 71691 32647 71733 32656
rect 71692 32562 71732 32647
rect 71499 32444 71541 32453
rect 71499 32404 71500 32444
rect 71540 32404 71541 32444
rect 71499 32395 71541 32404
rect 71595 32360 71637 32369
rect 71595 32320 71596 32360
rect 71636 32320 71637 32360
rect 71595 32311 71637 32320
rect 71596 32192 71636 32311
rect 71636 32152 71732 32192
rect 71596 32143 71636 32152
rect 71307 31352 71349 31361
rect 71307 31312 71308 31352
rect 71348 31312 71349 31352
rect 71307 31303 71349 31312
rect 71404 31352 71444 31361
rect 71211 30848 71253 30857
rect 71020 30808 71156 30848
rect 70924 30680 70964 30689
rect 70924 30185 70964 30640
rect 70923 30176 70965 30185
rect 70923 30136 70924 30176
rect 70964 30136 70965 30176
rect 70923 30127 70965 30136
rect 70828 29791 70868 29800
rect 71019 29840 71061 29849
rect 71019 29800 71020 29840
rect 71060 29800 71061 29840
rect 71019 29791 71061 29800
rect 71116 29840 71156 30808
rect 71211 30808 71212 30848
rect 71252 30808 71253 30848
rect 71211 30799 71253 30808
rect 71308 30773 71348 31303
rect 71307 30764 71349 30773
rect 71307 30724 71308 30764
rect 71348 30724 71349 30764
rect 71307 30715 71349 30724
rect 71212 30680 71252 30689
rect 71212 30437 71252 30640
rect 71308 30630 71348 30715
rect 71404 30521 71444 31312
rect 71596 31352 71636 31361
rect 71500 31268 71540 31277
rect 71403 30512 71445 30521
rect 71308 30472 71404 30512
rect 71444 30472 71445 30512
rect 71211 30428 71253 30437
rect 71211 30388 71212 30428
rect 71252 30388 71253 30428
rect 71211 30379 71253 30388
rect 71308 30260 71348 30472
rect 71403 30463 71445 30472
rect 71404 30378 71444 30463
rect 71500 30260 71540 31228
rect 71596 30512 71636 31312
rect 71596 30463 71636 30472
rect 71692 30269 71732 32152
rect 71788 30848 71828 33100
rect 71980 32864 72020 33412
rect 72076 33140 72116 33664
rect 72172 33655 72212 33664
rect 72268 33704 72308 33715
rect 72460 33713 72500 33798
rect 72268 33629 72308 33664
rect 72459 33704 72501 33713
rect 72459 33664 72460 33704
rect 72500 33664 72501 33704
rect 72459 33655 72501 33664
rect 72652 33704 72692 33713
rect 72267 33620 72309 33629
rect 72267 33580 72268 33620
rect 72308 33580 72309 33620
rect 72267 33571 72309 33580
rect 72555 33620 72597 33629
rect 72555 33580 72556 33620
rect 72596 33580 72597 33620
rect 72555 33571 72597 33580
rect 72556 33486 72596 33571
rect 72076 33100 72308 33140
rect 72172 32864 72212 32873
rect 71980 32824 72172 32864
rect 72172 32815 72212 32824
rect 71979 32696 72021 32705
rect 72268 32696 72308 33100
rect 72555 32864 72597 32873
rect 72555 32824 72556 32864
rect 72596 32824 72597 32864
rect 72555 32815 72597 32824
rect 72556 32730 72596 32815
rect 71979 32656 71980 32696
rect 72020 32656 72021 32696
rect 71979 32647 72021 32656
rect 72172 32656 72308 32696
rect 71883 32360 71925 32369
rect 71883 32320 71884 32360
rect 71924 32320 71925 32360
rect 71883 32311 71925 32320
rect 71884 32192 71924 32311
rect 71980 32276 72020 32647
rect 72075 32528 72117 32537
rect 72075 32488 72076 32528
rect 72116 32488 72117 32528
rect 72075 32479 72117 32488
rect 71980 32227 72020 32236
rect 71884 32143 71924 32152
rect 71788 30808 71924 30848
rect 71788 30680 71828 30689
rect 71116 29791 71156 29800
rect 71212 30220 71348 30260
rect 71404 30220 71540 30260
rect 71691 30260 71733 30269
rect 71691 30220 71692 30260
rect 71732 30220 71733 30260
rect 70923 29756 70965 29765
rect 70923 29716 70924 29756
rect 70964 29716 70965 29756
rect 70923 29707 70965 29716
rect 70924 29622 70964 29707
rect 71020 29706 71060 29791
rect 70923 29420 70965 29429
rect 70923 29380 70924 29420
rect 70964 29380 70965 29420
rect 70923 29371 70965 29380
rect 70732 29177 70772 29296
rect 70731 29168 70773 29177
rect 70731 29128 70732 29168
rect 70772 29128 70773 29168
rect 70731 29119 70773 29128
rect 70924 29084 70964 29371
rect 70924 29035 70964 29044
rect 71115 29084 71157 29093
rect 71115 29044 71116 29084
rect 71156 29044 71157 29084
rect 71115 29035 71157 29044
rect 71116 28950 71156 29035
rect 71212 28925 71252 30220
rect 71404 29849 71444 30220
rect 71691 30211 71733 30220
rect 71500 30092 71540 30101
rect 71788 30092 71828 30640
rect 71540 30052 71828 30092
rect 71500 30043 71540 30052
rect 71884 30008 71924 30808
rect 72076 30185 72116 32479
rect 72172 32033 72212 32656
rect 72652 32369 72692 33664
rect 72651 32360 72693 32369
rect 72651 32320 72652 32360
rect 72692 32320 72693 32360
rect 72651 32311 72693 32320
rect 72748 32201 72788 33916
rect 72844 33452 72884 36679
rect 72939 36476 72981 36485
rect 72939 36436 72940 36476
rect 72980 36436 72981 36476
rect 72939 36427 72981 36436
rect 72940 35720 72980 36427
rect 73035 35972 73077 35981
rect 73035 35932 73036 35972
rect 73076 35932 73077 35972
rect 73132 35972 73172 37948
rect 73611 37484 73653 37493
rect 73611 37444 73612 37484
rect 73652 37444 73748 37484
rect 73611 37435 73653 37444
rect 73227 37400 73269 37409
rect 73227 37360 73228 37400
rect 73268 37360 73269 37400
rect 73227 37351 73269 37360
rect 73420 37358 73460 37411
rect 73228 36905 73268 37351
rect 73419 37318 73420 37325
rect 73516 37400 73556 37409
rect 73460 37318 73461 37325
rect 73419 37316 73461 37318
rect 73419 37276 73420 37316
rect 73460 37276 73461 37316
rect 73419 37267 73461 37276
rect 73324 37232 73364 37241
rect 73324 36980 73364 37192
rect 73516 37064 73556 37360
rect 73708 37400 73748 37444
rect 73708 37351 73748 37360
rect 73900 37400 73940 37411
rect 73900 37325 73940 37360
rect 73995 37400 74037 37409
rect 73995 37360 73996 37400
rect 74036 37360 74037 37400
rect 73995 37351 74037 37360
rect 73899 37316 73941 37325
rect 73899 37276 73900 37316
rect 73940 37276 73941 37316
rect 73899 37267 73941 37276
rect 73996 37266 74036 37351
rect 73804 37232 73844 37241
rect 73516 37024 73748 37064
rect 73324 36940 73556 36980
rect 73227 36896 73269 36905
rect 73227 36856 73228 36896
rect 73268 36856 73269 36896
rect 73227 36847 73269 36856
rect 73323 36812 73365 36821
rect 73323 36772 73324 36812
rect 73364 36772 73365 36812
rect 73323 36763 73365 36772
rect 73516 36812 73556 36940
rect 73516 36763 73556 36772
rect 73324 36678 73364 36763
rect 73515 36560 73557 36569
rect 73515 36520 73516 36560
rect 73556 36520 73557 36560
rect 73515 36511 73557 36520
rect 73516 36065 73556 36511
rect 73708 36140 73748 37024
rect 73804 36821 73844 37192
rect 74092 37148 74132 38032
rect 75916 38032 76012 38072
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 73900 37108 74132 37148
rect 74284 37400 74324 37409
rect 73803 36812 73845 36821
rect 73803 36772 73804 36812
rect 73844 36772 73845 36812
rect 73803 36763 73845 36772
rect 73900 36728 73940 37108
rect 74091 36980 74133 36989
rect 74091 36940 74092 36980
rect 74132 36940 74133 36980
rect 74091 36931 74133 36940
rect 73900 36679 73940 36688
rect 73708 36091 73748 36100
rect 74092 36140 74132 36931
rect 74284 36149 74324 37360
rect 74476 37400 74516 37409
rect 74379 37316 74421 37325
rect 74379 37276 74380 37316
rect 74420 37276 74421 37316
rect 74379 37267 74421 37276
rect 74380 37182 74420 37267
rect 74476 36233 74516 37360
rect 74572 37400 74612 37409
rect 74572 37241 74612 37360
rect 74763 37400 74805 37409
rect 74763 37360 74764 37400
rect 74804 37360 74805 37400
rect 74763 37351 74805 37360
rect 75052 37400 75092 37409
rect 74571 37232 74613 37241
rect 74571 37192 74572 37232
rect 74612 37192 74613 37232
rect 74571 37183 74613 37192
rect 74764 36728 74804 37351
rect 75052 37241 75092 37360
rect 75148 37400 75188 37409
rect 75051 37232 75093 37241
rect 75051 37192 75052 37232
rect 75092 37192 75093 37232
rect 75051 37183 75093 37192
rect 75148 36737 75188 37360
rect 75244 37400 75284 37409
rect 75244 36905 75284 37360
rect 75916 37400 75956 38032
rect 76012 38023 76052 38032
rect 75916 37351 75956 37360
rect 76779 37400 76821 37409
rect 76779 37360 76780 37400
rect 76820 37360 76821 37400
rect 76779 37351 76821 37360
rect 75532 37316 75572 37325
rect 75572 37276 75860 37316
rect 75532 37267 75572 37276
rect 75340 37232 75380 37241
rect 75380 37192 75476 37232
rect 75340 37183 75380 37192
rect 75243 36896 75285 36905
rect 75243 36856 75244 36896
rect 75284 36856 75285 36896
rect 75243 36847 75285 36856
rect 74475 36224 74517 36233
rect 74475 36184 74476 36224
rect 74516 36184 74517 36224
rect 74475 36175 74517 36184
rect 74092 36091 74132 36100
rect 74283 36140 74325 36149
rect 74283 36100 74284 36140
rect 74324 36100 74325 36140
rect 74283 36091 74325 36100
rect 74764 36065 74804 36688
rect 75147 36728 75189 36737
rect 75147 36688 75148 36728
rect 75188 36688 75189 36728
rect 75147 36679 75189 36688
rect 75244 36569 75284 36847
rect 75436 36728 75476 37192
rect 75820 36980 75860 37276
rect 76780 37266 76820 37351
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 75820 36940 76244 36980
rect 76204 36896 76244 36940
rect 76204 36847 76244 36856
rect 76587 36812 76629 36821
rect 76587 36772 76588 36812
rect 76628 36772 76629 36812
rect 76587 36763 76629 36772
rect 76108 36728 76148 36737
rect 75436 36688 76108 36728
rect 76108 36679 76148 36688
rect 76203 36728 76245 36737
rect 76203 36688 76204 36728
rect 76244 36688 76245 36728
rect 76203 36679 76245 36688
rect 76300 36728 76340 36739
rect 75243 36560 75285 36569
rect 75243 36520 75244 36560
rect 75284 36520 75285 36560
rect 75243 36511 75285 36520
rect 76107 36560 76149 36569
rect 76107 36520 76108 36560
rect 76148 36520 76149 36560
rect 76107 36511 76149 36520
rect 75916 36476 75956 36485
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 73515 36056 73557 36065
rect 74668 36056 74708 36065
rect 73420 36014 73460 36023
rect 73515 36016 73516 36056
rect 73556 36016 73557 36056
rect 73515 36007 73557 36016
rect 74572 36016 74668 36056
rect 73132 35932 73364 35972
rect 73035 35923 73077 35932
rect 73036 35888 73076 35923
rect 73036 35837 73076 35848
rect 73132 35804 73172 35813
rect 73132 35720 73172 35764
rect 72940 35680 73172 35720
rect 73035 35300 73077 35309
rect 73035 35260 73036 35300
rect 73076 35260 73077 35300
rect 73035 35251 73077 35260
rect 72844 33412 72980 33452
rect 72843 32864 72885 32873
rect 72843 32824 72844 32864
rect 72884 32824 72885 32864
rect 72843 32815 72885 32824
rect 72460 32192 72500 32201
rect 72268 32152 72460 32192
rect 72171 32024 72213 32033
rect 72171 31984 72172 32024
rect 72212 31984 72213 32024
rect 72171 31975 72213 31984
rect 72268 32024 72308 32152
rect 72460 32143 72500 32152
rect 72652 32192 72692 32201
rect 72652 32117 72692 32152
rect 72747 32192 72789 32201
rect 72747 32152 72748 32192
rect 72788 32152 72789 32192
rect 72747 32143 72789 32152
rect 72651 32108 72693 32117
rect 72651 32068 72652 32108
rect 72692 32068 72693 32108
rect 72651 32059 72693 32068
rect 72268 31975 72308 31984
rect 72555 32024 72597 32033
rect 72555 31984 72556 32024
rect 72596 31984 72597 32024
rect 72555 31975 72597 31984
rect 72556 31890 72596 31975
rect 72363 31772 72405 31781
rect 72363 31732 72364 31772
rect 72404 31732 72405 31772
rect 72363 31723 72405 31732
rect 72268 31520 72308 31529
rect 72172 31480 72268 31520
rect 72172 30680 72212 31480
rect 72268 31471 72308 31480
rect 72172 30631 72212 30640
rect 72171 30428 72213 30437
rect 72171 30388 72172 30428
rect 72212 30388 72213 30428
rect 72171 30379 72213 30388
rect 72075 30176 72117 30185
rect 72075 30136 72076 30176
rect 72116 30136 72117 30176
rect 72075 30127 72117 30136
rect 71596 29968 71924 30008
rect 71403 29840 71445 29849
rect 71403 29800 71404 29840
rect 71444 29800 71445 29840
rect 71403 29791 71445 29800
rect 71500 29840 71540 29849
rect 71596 29840 71636 29968
rect 71540 29800 71636 29840
rect 71692 29840 71732 29849
rect 71500 29791 71540 29800
rect 71307 29756 71349 29765
rect 71307 29716 71308 29756
rect 71348 29716 71349 29756
rect 71307 29707 71349 29716
rect 71308 29009 71348 29707
rect 71404 29672 71444 29791
rect 71692 29672 71732 29800
rect 71787 29840 71829 29849
rect 71787 29800 71788 29840
rect 71828 29800 71829 29840
rect 71787 29791 71829 29800
rect 71788 29706 71828 29791
rect 71404 29632 71732 29672
rect 71884 29345 71924 29968
rect 71979 29924 72021 29933
rect 71979 29884 71980 29924
rect 72020 29884 72021 29924
rect 71979 29875 72021 29884
rect 71980 29840 72020 29875
rect 71980 29789 72020 29800
rect 72075 29840 72117 29849
rect 72075 29800 72076 29840
rect 72116 29800 72117 29840
rect 72075 29791 72117 29800
rect 72172 29840 72212 30379
rect 72267 30176 72309 30185
rect 72267 30136 72268 30176
rect 72308 30136 72309 30176
rect 72267 30127 72309 30136
rect 72172 29791 72212 29800
rect 72076 29706 72116 29791
rect 72268 29429 72308 30127
rect 72267 29420 72309 29429
rect 72267 29380 72268 29420
rect 72308 29380 72309 29420
rect 72267 29371 72309 29380
rect 71692 29336 71732 29345
rect 71883 29336 71925 29345
rect 71404 29296 71692 29336
rect 71732 29296 71884 29336
rect 71924 29296 71925 29336
rect 71307 29000 71349 29009
rect 71307 28960 71308 29000
rect 71348 28960 71349 29000
rect 71307 28951 71349 28960
rect 70827 28916 70869 28925
rect 70827 28876 70828 28916
rect 70868 28876 70869 28916
rect 70827 28867 70869 28876
rect 71211 28916 71253 28925
rect 71211 28876 71212 28916
rect 71252 28876 71253 28916
rect 71211 28867 71253 28876
rect 70636 28540 70772 28580
rect 70252 28279 70292 28288
rect 70348 28456 70676 28496
rect 69580 27868 70196 27908
rect 69483 27859 69525 27868
rect 69387 27824 69429 27833
rect 69387 27784 69388 27824
rect 69428 27784 69429 27824
rect 69387 27775 69429 27784
rect 69100 27700 69236 27740
rect 68907 27488 68949 27497
rect 68907 27448 68908 27488
rect 68948 27448 68949 27488
rect 68907 27439 68949 27448
rect 68811 27236 68853 27245
rect 68811 27196 68812 27236
rect 68852 27196 68853 27236
rect 68811 27187 68853 27196
rect 68812 27068 68852 27077
rect 68908 27068 68948 27439
rect 69003 27236 69045 27245
rect 69003 27196 69004 27236
rect 69044 27196 69045 27236
rect 69003 27187 69045 27196
rect 68852 27028 68948 27068
rect 68812 27019 68852 27028
rect 69004 26900 69044 27187
rect 69004 26851 69044 26860
rect 68907 26816 68949 26825
rect 68907 26776 68908 26816
rect 68948 26776 68949 26816
rect 68907 26767 68949 26776
rect 68811 26564 68853 26573
rect 68811 26524 68812 26564
rect 68852 26524 68853 26564
rect 68811 26515 68853 26524
rect 68812 26060 68852 26515
rect 68812 26011 68852 26020
rect 68908 23969 68948 26767
rect 69003 26312 69045 26321
rect 69003 26272 69004 26312
rect 69044 26272 69045 26312
rect 69003 26263 69045 26272
rect 68907 23960 68949 23969
rect 68812 23920 68908 23960
rect 68948 23920 68949 23960
rect 68524 23743 68564 23752
rect 68715 23792 68757 23801
rect 68715 23752 68716 23792
rect 68756 23752 68757 23792
rect 68715 23743 68757 23752
rect 68620 23624 68660 23633
rect 68620 23060 68660 23584
rect 68812 23060 68852 23920
rect 68907 23911 68949 23920
rect 68908 23792 68948 23801
rect 69004 23792 69044 26263
rect 68948 23752 69044 23792
rect 69100 23792 69140 27700
rect 69772 27665 69812 27750
rect 70059 27740 70101 27749
rect 70059 27700 70060 27740
rect 70100 27700 70101 27740
rect 70059 27691 70101 27700
rect 69580 27656 69620 27665
rect 69771 27656 69813 27665
rect 69196 27616 69524 27656
rect 69196 26816 69236 27616
rect 69388 27488 69428 27497
rect 69484 27488 69524 27616
rect 69620 27616 69716 27656
rect 69580 27607 69620 27616
rect 69580 27488 69620 27497
rect 69484 27448 69580 27488
rect 69388 26816 69428 27448
rect 69580 27439 69620 27448
rect 69580 26816 69620 26825
rect 69388 26776 69580 26816
rect 69196 26767 69236 26776
rect 69580 26767 69620 26776
rect 69387 26480 69429 26489
rect 69387 26440 69388 26480
rect 69428 26440 69429 26480
rect 69387 26431 69429 26440
rect 69291 26144 69333 26153
rect 69291 26104 69292 26144
rect 69332 26104 69333 26144
rect 69291 26095 69333 26104
rect 69388 26144 69428 26431
rect 69580 26312 69620 26321
rect 69676 26312 69716 27616
rect 69771 27616 69772 27656
rect 69812 27616 69813 27656
rect 69771 27607 69813 27616
rect 69868 27656 69908 27665
rect 69771 27488 69813 27497
rect 69771 27448 69772 27488
rect 69812 27448 69813 27488
rect 69868 27488 69908 27616
rect 70060 27656 70100 27691
rect 70060 27605 70100 27616
rect 70060 27488 70100 27497
rect 69868 27448 70060 27488
rect 69771 27439 69813 27448
rect 70060 27439 70100 27448
rect 69620 26272 69716 26312
rect 69580 26263 69620 26272
rect 69483 26228 69525 26237
rect 69483 26188 69484 26228
rect 69524 26188 69525 26228
rect 69483 26179 69525 26188
rect 69388 26095 69428 26104
rect 69484 26144 69524 26179
rect 69292 26010 69332 26095
rect 69484 26093 69524 26104
rect 69195 25304 69237 25313
rect 69195 25264 69196 25304
rect 69236 25264 69237 25304
rect 69195 25255 69237 25264
rect 69196 25170 69236 25255
rect 69292 23792 69332 23801
rect 69772 23792 69812 27439
rect 70156 23969 70196 27868
rect 70251 27740 70293 27749
rect 70251 27700 70252 27740
rect 70292 27700 70293 27740
rect 70251 27691 70293 27700
rect 70252 27656 70292 27691
rect 70252 27413 70292 27616
rect 70348 27656 70388 28456
rect 70539 28328 70581 28337
rect 70539 28288 70540 28328
rect 70580 28288 70581 28328
rect 70539 28279 70581 28288
rect 70636 28328 70676 28456
rect 70636 28279 70676 28288
rect 70540 28194 70580 28279
rect 70635 28160 70677 28169
rect 70635 28120 70636 28160
rect 70676 28120 70677 28160
rect 70635 28111 70677 28120
rect 70539 27908 70581 27917
rect 70539 27868 70540 27908
rect 70580 27868 70581 27908
rect 70539 27859 70581 27868
rect 70348 27607 70388 27616
rect 70251 27404 70293 27413
rect 70251 27364 70252 27404
rect 70292 27364 70293 27404
rect 70251 27355 70293 27364
rect 70444 26816 70484 26825
rect 70348 26776 70444 26816
rect 70348 25313 70388 26776
rect 70444 26767 70484 26776
rect 70443 26648 70485 26657
rect 70443 26608 70444 26648
rect 70484 26608 70485 26648
rect 70443 26599 70485 26608
rect 70444 26060 70484 26599
rect 70444 26011 70484 26020
rect 70540 26312 70580 27859
rect 70636 27656 70676 28111
rect 70636 27607 70676 27616
rect 70732 27740 70772 28540
rect 70828 28169 70868 28867
rect 71308 28866 71348 28951
rect 71404 28748 71444 29296
rect 71692 29287 71732 29296
rect 71883 29287 71925 29296
rect 71884 29202 71924 29287
rect 71499 29168 71541 29177
rect 72364 29168 72404 31723
rect 72652 30521 72692 32059
rect 72844 32024 72884 32815
rect 72940 32537 72980 33412
rect 72939 32528 72981 32537
rect 72939 32488 72940 32528
rect 72980 32488 72981 32528
rect 72939 32479 72981 32488
rect 72939 32360 72981 32369
rect 72939 32320 72940 32360
rect 72980 32320 72981 32360
rect 72939 32311 72981 32320
rect 72844 31975 72884 31984
rect 72940 31865 72980 32311
rect 73036 32117 73076 35251
rect 73227 35132 73269 35141
rect 73227 35092 73228 35132
rect 73268 35092 73269 35132
rect 73227 35083 73269 35092
rect 73131 32948 73173 32957
rect 73131 32908 73132 32948
rect 73172 32908 73173 32948
rect 73131 32899 73173 32908
rect 73035 32108 73077 32117
rect 73035 32068 73036 32108
rect 73076 32068 73077 32108
rect 73035 32059 73077 32068
rect 72939 31856 72981 31865
rect 72939 31816 72940 31856
rect 72980 31816 72981 31856
rect 72939 31807 72981 31816
rect 73035 31688 73077 31697
rect 73035 31648 73036 31688
rect 73076 31648 73077 31688
rect 73035 31639 73077 31648
rect 73036 31361 73076 31639
rect 73035 31352 73077 31361
rect 73035 31312 73036 31352
rect 73076 31312 73077 31352
rect 73035 31303 73077 31312
rect 73036 30680 73076 31303
rect 73036 30631 73076 30640
rect 72651 30512 72693 30521
rect 72651 30472 72652 30512
rect 72692 30472 72693 30512
rect 72651 30463 72693 30472
rect 72459 30260 72501 30269
rect 72459 30220 72460 30260
rect 72500 30220 72501 30260
rect 72459 30211 72501 30220
rect 72460 29177 72500 30211
rect 72555 29420 72597 29429
rect 72555 29380 72556 29420
rect 72596 29380 72597 29420
rect 72555 29371 72597 29380
rect 71499 29128 71500 29168
rect 71540 29128 71541 29168
rect 71499 29119 71541 29128
rect 72076 29128 72404 29168
rect 72459 29168 72501 29177
rect 72459 29128 72460 29168
rect 72500 29128 72501 29168
rect 71020 28708 71444 28748
rect 71500 29084 71540 29119
rect 70924 28496 70964 28505
rect 70827 28160 70869 28169
rect 70827 28120 70828 28160
rect 70868 28120 70869 28160
rect 70827 28111 70869 28120
rect 70732 27488 70772 27700
rect 70828 27656 70868 27665
rect 70924 27656 70964 28456
rect 70868 27616 70964 27656
rect 71020 27656 71060 28708
rect 71404 28244 71444 28253
rect 71116 27824 71156 27833
rect 71404 27824 71444 28204
rect 71500 27917 71540 29044
rect 71979 29084 72021 29093
rect 71979 29044 71980 29084
rect 72020 29044 72021 29084
rect 71979 29035 72021 29044
rect 72076 29084 72116 29128
rect 72076 29035 72116 29044
rect 71883 28916 71925 28925
rect 71883 28876 71884 28916
rect 71924 28876 71925 28916
rect 71883 28867 71925 28876
rect 71884 28782 71924 28867
rect 71691 28412 71733 28421
rect 71691 28372 71692 28412
rect 71732 28372 71733 28412
rect 71691 28363 71733 28372
rect 71499 27908 71541 27917
rect 71499 27868 71500 27908
rect 71540 27868 71541 27908
rect 71499 27859 71541 27868
rect 71156 27784 71444 27824
rect 71116 27775 71156 27784
rect 71500 27749 71540 27780
rect 71499 27740 71541 27749
rect 71499 27700 71500 27740
rect 71540 27700 71541 27740
rect 71499 27691 71541 27700
rect 70828 27607 70868 27616
rect 71020 27607 71060 27616
rect 71212 27656 71252 27665
rect 71212 27488 71252 27616
rect 70732 27448 71252 27488
rect 71308 27656 71348 27665
rect 71308 27413 71348 27616
rect 71500 27656 71540 27691
rect 71692 27669 71732 28363
rect 71788 28328 71828 28337
rect 71828 28288 71924 28328
rect 71788 28279 71828 28288
rect 71692 27620 71732 27629
rect 71787 27656 71829 27665
rect 71307 27404 71349 27413
rect 71307 27364 71308 27404
rect 71348 27364 71349 27404
rect 71307 27355 71349 27364
rect 70827 27320 70869 27329
rect 70827 27280 70828 27320
rect 70868 27280 70869 27320
rect 70827 27271 70869 27280
rect 71403 27320 71445 27329
rect 71403 27280 71404 27320
rect 71444 27280 71445 27320
rect 71403 27271 71445 27280
rect 70636 26312 70676 26321
rect 70540 26272 70636 26312
rect 70347 25304 70389 25313
rect 70347 25264 70348 25304
rect 70388 25264 70389 25304
rect 70347 25255 70389 25264
rect 70347 25136 70389 25145
rect 70347 25096 70348 25136
rect 70388 25096 70389 25136
rect 70347 25087 70389 25096
rect 70348 24809 70388 25087
rect 70540 24893 70580 26272
rect 70636 26263 70676 26272
rect 70828 25976 70868 27271
rect 70923 26648 70965 26657
rect 70923 26608 70924 26648
rect 70964 26608 70965 26648
rect 70923 26599 70965 26608
rect 70924 26144 70964 26599
rect 71307 26312 71349 26321
rect 71307 26272 71308 26312
rect 71348 26272 71349 26312
rect 71307 26263 71349 26272
rect 71308 26228 71348 26263
rect 71308 26153 71348 26188
rect 70924 26095 70964 26104
rect 71212 26144 71252 26153
rect 70828 25936 70964 25976
rect 70636 25220 70676 25229
rect 70539 24884 70581 24893
rect 70539 24844 70540 24884
rect 70580 24844 70581 24884
rect 70539 24835 70581 24844
rect 70347 24800 70389 24809
rect 70347 24760 70348 24800
rect 70388 24760 70389 24800
rect 70347 24751 70389 24760
rect 70540 24632 70580 24835
rect 70636 24800 70676 25180
rect 70828 24800 70868 24809
rect 70636 24760 70828 24800
rect 70828 24751 70868 24760
rect 70732 24632 70772 24641
rect 70540 24592 70732 24632
rect 70732 24583 70772 24592
rect 70924 24632 70964 25936
rect 71212 25481 71252 26104
rect 71307 26144 71349 26153
rect 71307 26104 71308 26144
rect 71348 26104 71349 26144
rect 71307 26095 71349 26104
rect 71308 26064 71348 26095
rect 71211 25472 71253 25481
rect 71211 25432 71212 25472
rect 71252 25432 71253 25472
rect 71211 25423 71253 25432
rect 71020 25304 71060 25313
rect 71060 25264 71252 25304
rect 71020 25255 71060 25264
rect 70924 24583 70964 24592
rect 71019 24632 71061 24641
rect 71019 24592 71020 24632
rect 71060 24592 71061 24632
rect 71019 24583 71061 24592
rect 71020 24498 71060 24583
rect 71212 24464 71252 25264
rect 71212 24415 71252 24424
rect 70155 23960 70197 23969
rect 70155 23920 70156 23960
rect 70196 23920 70197 23960
rect 70155 23911 70197 23920
rect 70539 23960 70581 23969
rect 70539 23920 70540 23960
rect 70580 23920 70581 23960
rect 70539 23911 70581 23920
rect 70827 23960 70869 23969
rect 70827 23920 70828 23960
rect 70868 23920 70869 23960
rect 70827 23911 70869 23920
rect 70155 23792 70197 23801
rect 69100 23752 69292 23792
rect 69332 23752 69620 23792
rect 68908 23633 68948 23752
rect 69292 23743 69332 23752
rect 68907 23624 68949 23633
rect 68907 23584 68908 23624
rect 68948 23584 68949 23624
rect 68907 23575 68949 23584
rect 69004 23624 69044 23633
rect 69004 23060 69044 23584
rect 69291 23624 69333 23633
rect 69291 23584 69292 23624
rect 69332 23584 69333 23624
rect 69291 23575 69333 23584
rect 69388 23624 69428 23633
rect 69292 23060 69332 23575
rect 68044 23020 68095 23060
rect 68236 23020 68385 23060
rect 68428 23020 68495 23060
rect 68620 23020 68756 23060
rect 68812 23020 68895 23060
rect 69004 23020 69185 23060
rect 67852 22744 67985 22784
rect 67655 22596 67695 22744
rect 67945 22596 67985 22744
rect 68055 22596 68095 23020
rect 68345 22596 68385 23020
rect 68455 22596 68495 23020
rect 68716 22784 68756 23020
rect 68716 22744 68785 22784
rect 68745 22596 68785 22744
rect 68855 22596 68895 23020
rect 69145 22596 69185 23020
rect 69255 23020 69332 23060
rect 69388 23060 69428 23584
rect 69580 23060 69620 23752
rect 69812 23752 70100 23792
rect 69772 23743 69812 23752
rect 69868 23624 69908 23633
rect 69868 23060 69908 23584
rect 70060 23060 70100 23752
rect 70155 23752 70156 23792
rect 70196 23752 70197 23792
rect 70155 23743 70197 23752
rect 70443 23792 70485 23801
rect 70443 23752 70444 23792
rect 70484 23752 70485 23792
rect 70443 23743 70485 23752
rect 70540 23792 70580 23911
rect 70540 23743 70580 23752
rect 70156 23658 70196 23743
rect 69388 23020 69524 23060
rect 69580 23020 69695 23060
rect 69868 23020 69985 23060
rect 69255 22596 69295 23020
rect 69484 22784 69524 23020
rect 69484 22744 69585 22784
rect 69545 22596 69585 22744
rect 69655 22596 69695 23020
rect 69945 22596 69985 23020
rect 70055 23020 70100 23060
rect 70252 23624 70292 23633
rect 70252 23060 70292 23584
rect 70444 23060 70484 23743
rect 70636 23624 70676 23633
rect 70636 23060 70676 23584
rect 70828 23060 70868 23911
rect 70923 23792 70965 23801
rect 71308 23792 71348 23801
rect 71404 23792 71444 27271
rect 71500 24800 71540 27616
rect 71787 27616 71788 27656
rect 71828 27616 71829 27656
rect 71787 27607 71829 27616
rect 71595 27404 71637 27413
rect 71595 27364 71596 27404
rect 71636 27364 71637 27404
rect 71595 27355 71637 27364
rect 71596 27270 71636 27355
rect 71788 27068 71828 27607
rect 71884 27488 71924 28288
rect 71884 27439 71924 27448
rect 71980 27068 72020 29035
rect 71788 27028 71924 27068
rect 71788 26900 71828 26909
rect 71596 26648 71636 26657
rect 71596 26321 71636 26608
rect 71788 26321 71828 26860
rect 71595 26312 71637 26321
rect 71595 26272 71596 26312
rect 71636 26272 71637 26312
rect 71595 26263 71637 26272
rect 71787 26312 71829 26321
rect 71787 26272 71788 26312
rect 71828 26272 71829 26312
rect 71787 26263 71829 26272
rect 71884 26228 71924 27028
rect 71980 27019 72020 27028
rect 72172 27068 72212 29128
rect 72459 29119 72501 29128
rect 72172 27019 72212 27028
rect 72364 26900 72404 26909
rect 72364 26741 72404 26860
rect 72363 26732 72405 26741
rect 72363 26692 72364 26732
rect 72404 26692 72405 26732
rect 72363 26683 72405 26692
rect 71979 26648 72021 26657
rect 72172 26648 72212 26657
rect 71979 26608 71980 26648
rect 72020 26608 72021 26648
rect 71979 26599 72021 26608
rect 72076 26608 72172 26648
rect 71980 26514 72020 26599
rect 72076 26396 72116 26608
rect 72172 26599 72212 26608
rect 72556 26489 72596 29371
rect 72652 28328 72692 28337
rect 72555 26480 72597 26489
rect 72555 26440 72556 26480
rect 72596 26440 72597 26480
rect 72555 26431 72597 26440
rect 71884 26179 71924 26188
rect 71980 26356 72116 26396
rect 71980 26153 72020 26356
rect 72556 26237 72596 26431
rect 72555 26228 72597 26237
rect 72555 26188 72556 26228
rect 72596 26188 72597 26228
rect 72555 26179 72597 26188
rect 71788 26144 71828 26153
rect 71596 25892 71636 25901
rect 71788 25892 71828 26104
rect 71979 26144 72021 26153
rect 71979 26104 71980 26144
rect 72020 26104 72021 26144
rect 71979 26095 72021 26104
rect 72652 25901 72692 28288
rect 73035 26900 73077 26909
rect 73035 26860 73036 26900
rect 73076 26860 73077 26900
rect 73035 26851 73077 26860
rect 73036 26816 73076 26851
rect 73036 26765 73076 26776
rect 71636 25852 71828 25892
rect 72651 25892 72693 25901
rect 72651 25852 72652 25892
rect 72692 25852 72693 25892
rect 71596 25843 71636 25852
rect 72651 25843 72693 25852
rect 71787 25472 71829 25481
rect 71787 25432 71788 25472
rect 71828 25432 71829 25472
rect 71787 25423 71829 25432
rect 71595 24800 71637 24809
rect 71500 24760 71596 24800
rect 71636 24760 71637 24800
rect 71595 24751 71637 24760
rect 71596 24632 71636 24751
rect 71596 24583 71636 24592
rect 71691 24632 71733 24641
rect 71691 24592 71692 24632
rect 71732 24592 71733 24632
rect 71691 24583 71733 24592
rect 71788 24632 71828 25423
rect 72652 25313 72692 25843
rect 72843 25472 72885 25481
rect 72843 25432 72844 25472
rect 72884 25432 72885 25472
rect 72843 25423 72885 25432
rect 73035 25472 73077 25481
rect 73035 25432 73036 25472
rect 73076 25432 73077 25472
rect 73035 25423 73077 25432
rect 71883 25304 71925 25313
rect 71883 25264 71884 25304
rect 71924 25264 71925 25304
rect 71883 25255 71925 25264
rect 72651 25304 72693 25313
rect 72651 25264 72652 25304
rect 72692 25264 72693 25304
rect 72651 25255 72693 25264
rect 71884 25170 71924 25255
rect 72459 25136 72501 25145
rect 72459 25096 72460 25136
rect 72500 25096 72501 25136
rect 72459 25087 72501 25096
rect 72075 24968 72117 24977
rect 72075 24928 72076 24968
rect 72116 24928 72117 24968
rect 72075 24919 72117 24928
rect 71788 24583 71828 24592
rect 71692 24498 71732 24583
rect 71691 23792 71733 23801
rect 70923 23752 70924 23792
rect 70964 23752 71252 23792
rect 70923 23743 70965 23752
rect 70924 23658 70964 23743
rect 71020 23624 71060 23633
rect 71020 23060 71060 23584
rect 71212 23060 71252 23752
rect 71348 23752 71636 23792
rect 71308 23743 71348 23752
rect 71404 23624 71444 23633
rect 71404 23060 71444 23584
rect 71596 23060 71636 23752
rect 71691 23752 71692 23792
rect 71732 23752 71733 23792
rect 71691 23743 71733 23752
rect 71979 23792 72021 23801
rect 71979 23752 71980 23792
rect 72020 23752 72021 23792
rect 71979 23743 72021 23752
rect 72076 23792 72116 24919
rect 72460 23792 72500 25087
rect 72844 23792 72884 25423
rect 73036 25338 73076 25423
rect 73132 24221 73172 32899
rect 73228 29093 73268 35083
rect 73324 33140 73364 35932
rect 73420 35897 73460 35974
rect 73419 35888 73461 35897
rect 73419 35848 73420 35888
rect 73460 35848 73461 35888
rect 73419 35839 73461 35848
rect 73516 35720 73556 36007
rect 73803 35972 73845 35981
rect 73803 35932 73804 35972
rect 73844 35932 73845 35972
rect 73803 35923 73845 35932
rect 73612 35888 73652 35897
rect 73804 35888 73844 35923
rect 73652 35848 73748 35888
rect 73612 35839 73652 35848
rect 73516 35680 73652 35720
rect 73453 34376 73493 34385
rect 73612 34376 73652 35680
rect 73708 35477 73748 35848
rect 73804 35837 73844 35848
rect 73995 35888 74037 35897
rect 73995 35848 73996 35888
rect 74036 35848 74037 35888
rect 73995 35839 74037 35848
rect 74188 35888 74228 35897
rect 74228 35848 74324 35888
rect 74188 35839 74228 35848
rect 73996 35754 74036 35839
rect 74284 35645 74324 35848
rect 74283 35636 74325 35645
rect 74283 35596 74284 35636
rect 74324 35596 74325 35636
rect 74283 35587 74325 35596
rect 73707 35468 73749 35477
rect 73707 35428 73708 35468
rect 73748 35428 73749 35468
rect 73707 35419 73749 35428
rect 74187 35216 74229 35225
rect 74187 35176 74188 35216
rect 74228 35176 74229 35216
rect 74187 35167 74229 35176
rect 74188 35082 74228 35167
rect 73493 34336 73652 34376
rect 73453 34327 73493 34336
rect 73707 33956 73749 33965
rect 73707 33916 73708 33956
rect 73748 33916 73749 33956
rect 73707 33907 73749 33916
rect 73708 33140 73748 33907
rect 73324 33100 73460 33140
rect 73708 33100 73844 33140
rect 73420 32853 73460 33100
rect 73420 32528 73460 32813
rect 73324 32488 73460 32528
rect 73324 31697 73364 32488
rect 73323 31688 73365 31697
rect 73323 31648 73324 31688
rect 73364 31648 73365 31688
rect 73323 31639 73365 31648
rect 73612 31268 73652 31277
rect 73515 31100 73557 31109
rect 73515 31060 73516 31100
rect 73556 31060 73557 31100
rect 73515 31051 73557 31060
rect 73420 29126 73460 29135
rect 73227 29084 73269 29093
rect 73227 29044 73228 29084
rect 73268 29044 73269 29084
rect 73227 29035 73269 29044
rect 73420 28589 73460 29086
rect 73419 28580 73461 28589
rect 73419 28540 73420 28580
rect 73460 28540 73461 28580
rect 73419 28531 73461 28540
rect 73516 27665 73556 31051
rect 73612 30857 73652 31228
rect 73611 30848 73653 30857
rect 73611 30808 73612 30848
rect 73652 30808 73653 30848
rect 73611 30799 73653 30808
rect 73707 30428 73749 30437
rect 73707 30388 73708 30428
rect 73748 30388 73749 30428
rect 73707 30379 73749 30388
rect 73515 27656 73557 27665
rect 73515 27616 73516 27656
rect 73556 27616 73557 27656
rect 73515 27607 73557 27616
rect 73516 27488 73556 27497
rect 73516 27152 73556 27448
rect 73420 27112 73556 27152
rect 73420 26852 73460 27112
rect 73420 26803 73460 26812
rect 73227 25976 73269 25985
rect 73227 25936 73228 25976
rect 73268 25936 73269 25976
rect 73227 25927 73269 25936
rect 73420 25934 73460 25943
rect 73228 25304 73268 25927
rect 73420 25640 73460 25894
rect 73420 25600 73556 25640
rect 73516 25304 73556 25600
rect 73612 25304 73652 25313
rect 73516 25264 73612 25304
rect 73228 25255 73268 25264
rect 73612 25255 73652 25264
rect 73131 24212 73173 24221
rect 73131 24172 73132 24212
rect 73172 24172 73173 24212
rect 73131 24163 73173 24172
rect 73323 23960 73365 23969
rect 73323 23920 73324 23960
rect 73364 23920 73365 23960
rect 73323 23911 73365 23920
rect 73611 23960 73653 23969
rect 73611 23920 73612 23960
rect 73652 23920 73653 23960
rect 73611 23911 73653 23920
rect 73324 23792 73364 23911
rect 72116 23752 72404 23792
rect 72076 23743 72116 23752
rect 71692 23658 71732 23743
rect 71788 23624 71828 23633
rect 71788 23060 71828 23584
rect 70252 23020 70385 23060
rect 70444 23020 70495 23060
rect 70636 23020 70785 23060
rect 70828 23020 70895 23060
rect 71020 23020 71156 23060
rect 71212 23020 71295 23060
rect 71404 23020 71540 23060
rect 71596 23020 71695 23060
rect 71788 23020 71924 23060
rect 70055 22596 70095 23020
rect 70345 22596 70385 23020
rect 70455 22596 70495 23020
rect 70745 22596 70785 23020
rect 70855 22596 70895 23020
rect 71116 22784 71156 23020
rect 71116 22744 71185 22784
rect 71145 22596 71185 22744
rect 71255 22596 71295 23020
rect 71500 22784 71540 23020
rect 71500 22744 71585 22784
rect 71545 22596 71585 22744
rect 71655 22596 71695 23020
rect 71884 22784 71924 23020
rect 71980 22868 72020 23743
rect 72172 23624 72212 23633
rect 72172 23060 72212 23584
rect 72364 23060 72404 23752
rect 72500 23752 72692 23792
rect 72460 23743 72500 23752
rect 72556 23624 72596 23633
rect 72172 23020 72308 23060
rect 72364 23020 72495 23060
rect 71980 22828 72116 22868
rect 72076 22784 72116 22828
rect 71884 22744 71985 22784
rect 71945 22596 71985 22744
rect 72055 22744 72116 22784
rect 72268 22784 72308 23020
rect 72268 22744 72385 22784
rect 72055 22596 72095 22744
rect 72345 22596 72385 22744
rect 72455 22596 72495 23020
rect 72556 22784 72596 23584
rect 72652 23060 72692 23752
rect 72884 23752 73268 23792
rect 72844 23743 72884 23752
rect 72940 23624 72980 23633
rect 72940 23060 72980 23584
rect 73228 23060 73268 23752
rect 73324 23743 73364 23752
rect 73420 23624 73460 23633
rect 73460 23584 73556 23624
rect 73420 23556 73460 23584
rect 72652 23020 72895 23060
rect 72940 23020 73185 23060
rect 73228 23020 73295 23060
rect 72556 22744 72785 22784
rect 72745 22596 72785 22744
rect 72855 22596 72895 23020
rect 73145 22596 73185 23020
rect 73255 22596 73295 23020
rect 73516 22784 73556 23584
rect 73612 23060 73652 23911
rect 73708 23792 73748 30379
rect 73804 30176 73844 33100
rect 74092 32024 74132 32033
rect 73996 31984 74092 32024
rect 73996 31352 74036 31984
rect 74092 31975 74132 31984
rect 74284 31781 74324 35587
rect 74572 35216 74612 36016
rect 74668 36007 74708 36016
rect 74763 36056 74805 36065
rect 74763 36016 74764 36056
rect 74804 36016 74805 36056
rect 74763 36007 74805 36016
rect 75435 36056 75477 36065
rect 75435 36016 75436 36056
rect 75476 36016 75477 36056
rect 75435 36007 75477 36016
rect 74572 35167 74612 35176
rect 75436 35216 75476 36007
rect 75916 35981 75956 36436
rect 75915 35972 75957 35981
rect 75915 35932 75916 35972
rect 75956 35932 75957 35972
rect 75915 35923 75957 35932
rect 75436 35167 75476 35176
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 74571 34208 74613 34217
rect 74571 34168 74572 34208
rect 74612 34168 74613 34208
rect 74571 34159 74613 34168
rect 75627 34208 75669 34217
rect 75627 34168 75628 34208
rect 75668 34168 75669 34208
rect 75627 34159 75669 34168
rect 74572 34074 74612 34159
rect 74859 33704 74901 33713
rect 74859 33664 74860 33704
rect 74900 33664 74901 33704
rect 74859 33655 74901 33664
rect 74763 33452 74805 33461
rect 74763 33412 74764 33452
rect 74804 33412 74805 33452
rect 74763 33403 74805 33412
rect 74764 32864 74804 33403
rect 74860 33209 74900 33655
rect 75052 33536 75092 33545
rect 74956 33496 75052 33536
rect 74859 33200 74901 33209
rect 74859 33160 74860 33200
rect 74900 33160 74901 33200
rect 74859 33151 74901 33160
rect 74764 32815 74804 32824
rect 74572 32696 74612 32705
rect 74572 31865 74612 32656
rect 74571 31856 74613 31865
rect 74571 31816 74572 31856
rect 74612 31816 74613 31856
rect 74860 31856 74900 33151
rect 74956 33140 74996 33496
rect 75052 33487 75092 33496
rect 75531 33536 75573 33545
rect 75531 33496 75532 33536
rect 75572 33496 75573 33536
rect 75531 33487 75573 33496
rect 75112 33284 75480 33293
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75112 33235 75480 33244
rect 74956 33100 75188 33140
rect 75148 32864 75188 33100
rect 75148 32815 75188 32824
rect 74860 31816 74996 31856
rect 74571 31807 74613 31816
rect 74283 31772 74325 31781
rect 74283 31732 74284 31772
rect 74324 31732 74325 31772
rect 74283 31723 74325 31732
rect 73996 31303 74036 31312
rect 74187 30428 74229 30437
rect 74187 30388 74188 30428
rect 74228 30388 74229 30428
rect 74187 30379 74229 30388
rect 74188 30294 74228 30379
rect 73804 30136 74036 30176
rect 73900 30008 73940 30017
rect 73804 29168 73844 29177
rect 73900 29168 73940 29968
rect 73844 29128 73940 29168
rect 73804 29119 73844 29128
rect 73803 28412 73845 28421
rect 73803 28372 73804 28412
rect 73844 28372 73845 28412
rect 73803 28363 73845 28372
rect 73804 23969 73844 28363
rect 73899 27656 73941 27665
rect 73899 27616 73900 27656
rect 73940 27616 73941 27656
rect 73899 27607 73941 27616
rect 73900 24053 73940 27607
rect 73899 24044 73941 24053
rect 73899 24004 73900 24044
rect 73940 24004 73941 24044
rect 73899 23995 73941 24004
rect 73996 23969 74036 30136
rect 74091 27404 74133 27413
rect 74091 27364 74092 27404
rect 74132 27364 74133 27404
rect 74091 27355 74133 27364
rect 74092 24632 74132 27355
rect 74284 26816 74324 26825
rect 74324 26776 74420 26816
rect 74284 26767 74324 26776
rect 74188 26144 74228 26153
rect 74188 24800 74228 26104
rect 74283 26144 74325 26153
rect 74283 26104 74284 26144
rect 74324 26104 74325 26144
rect 74283 26095 74325 26104
rect 74284 26010 74324 26095
rect 74380 25901 74420 26776
rect 74475 26312 74517 26321
rect 74475 26272 74476 26312
rect 74516 26272 74517 26312
rect 74475 26263 74517 26272
rect 74476 26144 74516 26263
rect 74476 26095 74516 26104
rect 74475 25976 74517 25985
rect 74475 25936 74476 25976
rect 74516 25936 74517 25976
rect 74475 25927 74517 25936
rect 74379 25892 74421 25901
rect 74379 25852 74380 25892
rect 74420 25852 74421 25892
rect 74379 25843 74421 25852
rect 74380 25304 74420 25843
rect 74476 25842 74516 25927
rect 74572 25388 74612 31807
rect 74859 31688 74901 31697
rect 74859 31648 74860 31688
rect 74900 31648 74901 31688
rect 74859 31639 74901 31648
rect 74667 31352 74709 31361
rect 74860 31352 74900 31639
rect 74667 31312 74668 31352
rect 74708 31312 74860 31352
rect 74667 31303 74709 31312
rect 74860 31303 74900 31312
rect 74668 29168 74708 31303
rect 74859 30764 74901 30773
rect 74859 30724 74860 30764
rect 74900 30724 74901 30764
rect 74859 30715 74901 30724
rect 74860 30630 74900 30715
rect 74956 30680 74996 31816
rect 75112 31772 75480 31781
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75112 31723 75480 31732
rect 75532 31100 75572 33487
rect 75244 31060 75572 31100
rect 75244 30932 75284 31060
rect 74956 30092 74996 30640
rect 75052 30892 75284 30932
rect 75052 30680 75092 30892
rect 75435 30848 75477 30857
rect 75435 30808 75436 30848
rect 75476 30808 75477 30848
rect 75628 30848 75668 34159
rect 75724 33704 75764 33713
rect 75724 32360 75764 33664
rect 75820 33704 75860 33715
rect 75820 33629 75860 33664
rect 75819 33620 75861 33629
rect 75819 33580 75820 33620
rect 75860 33580 75861 33620
rect 75819 33571 75861 33580
rect 75916 32528 75956 35923
rect 76108 35888 76148 36511
rect 76108 35839 76148 35848
rect 76204 35888 76244 36679
rect 76300 36653 76340 36688
rect 76396 36728 76436 36737
rect 76299 36644 76341 36653
rect 76299 36604 76300 36644
rect 76340 36604 76341 36644
rect 76299 36595 76341 36604
rect 76396 36140 76436 36688
rect 76588 36728 76628 36763
rect 76588 36677 76628 36688
rect 76780 36728 76820 36737
rect 76780 36653 76820 36688
rect 76875 36728 76917 36737
rect 76875 36688 76876 36728
rect 76916 36688 76917 36728
rect 76875 36679 76917 36688
rect 76779 36644 76821 36653
rect 76779 36604 76780 36644
rect 76820 36604 76821 36644
rect 76779 36595 76821 36604
rect 76587 36560 76629 36569
rect 76587 36520 76588 36560
rect 76628 36520 76629 36560
rect 76587 36511 76629 36520
rect 76588 36426 76628 36511
rect 76683 36224 76725 36233
rect 76683 36184 76684 36224
rect 76724 36184 76725 36224
rect 76683 36175 76725 36184
rect 76492 36140 76532 36149
rect 76396 36100 76492 36140
rect 76492 36091 76532 36100
rect 76492 35897 76532 35982
rect 76204 35839 76244 35848
rect 76300 35888 76340 35897
rect 76012 35720 76052 35729
rect 76300 35720 76340 35848
rect 76491 35888 76533 35897
rect 76491 35848 76492 35888
rect 76532 35848 76533 35888
rect 76491 35839 76533 35848
rect 76684 35888 76724 36175
rect 76780 36149 76820 36595
rect 76876 36594 76916 36679
rect 76779 36140 76821 36149
rect 76779 36100 76780 36140
rect 76820 36100 76821 36140
rect 76779 36091 76821 36100
rect 76972 36056 77012 38200
rect 77164 37409 77204 38200
rect 77260 38240 77300 38249
rect 77163 37400 77205 37409
rect 77163 37360 77164 37400
rect 77204 37360 77205 37400
rect 77163 37351 77205 37360
rect 77260 37241 77300 38200
rect 77548 37988 77588 37997
rect 77588 37948 77684 37988
rect 77548 37939 77588 37948
rect 77451 37400 77493 37409
rect 77451 37360 77452 37400
rect 77492 37360 77493 37400
rect 77451 37351 77493 37360
rect 77259 37232 77301 37241
rect 77259 37192 77260 37232
rect 77300 37192 77301 37232
rect 77259 37183 77301 37192
rect 77355 36812 77397 36821
rect 77355 36772 77356 36812
rect 77396 36772 77397 36812
rect 77355 36763 77397 36772
rect 77068 36728 77108 36737
rect 77068 36569 77108 36688
rect 77067 36560 77109 36569
rect 77067 36520 77068 36560
rect 77108 36520 77109 36560
rect 77067 36511 77109 36520
rect 76876 36016 77012 36056
rect 76684 35839 76724 35848
rect 76780 35888 76820 35897
rect 76780 35720 76820 35848
rect 76300 35680 76820 35720
rect 76012 34376 76052 35680
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 76107 35216 76149 35225
rect 76107 35176 76108 35216
rect 76148 35176 76149 35216
rect 76107 35167 76149 35176
rect 76012 34327 76052 34336
rect 76108 34292 76148 35167
rect 76491 35048 76533 35057
rect 76491 35008 76492 35048
rect 76532 35008 76533 35048
rect 76491 34999 76533 35008
rect 76492 34796 76532 34999
rect 76588 34964 76628 34973
rect 76588 34880 76628 34924
rect 76780 34880 76820 35680
rect 76876 35057 76916 36016
rect 77068 35888 77108 35897
rect 77068 35645 77108 35848
rect 77260 35888 77300 35897
rect 77164 35804 77204 35813
rect 77067 35636 77109 35645
rect 77067 35596 77068 35636
rect 77108 35596 77109 35636
rect 77067 35587 77109 35596
rect 77164 35393 77204 35764
rect 77163 35384 77205 35393
rect 77163 35344 77164 35384
rect 77204 35344 77205 35384
rect 77163 35335 77205 35344
rect 77068 35216 77108 35225
rect 77108 35176 77204 35216
rect 77068 35167 77108 35176
rect 76875 35048 76917 35057
rect 76875 35008 76876 35048
rect 76916 35008 76917 35048
rect 76875 34999 76917 35008
rect 76588 34840 77012 34880
rect 76492 34756 76628 34796
rect 76203 34376 76245 34385
rect 76203 34336 76204 34376
rect 76244 34336 76245 34376
rect 76203 34327 76245 34336
rect 76300 34376 76340 34385
rect 76588 34376 76628 34756
rect 76340 34336 76532 34376
rect 76300 34327 76340 34336
rect 76108 34243 76148 34252
rect 76204 34242 76244 34327
rect 76492 34208 76532 34336
rect 76588 34327 76628 34336
rect 76876 34376 76916 34387
rect 76876 34301 76916 34336
rect 76972 34376 77012 34840
rect 77164 34460 77204 35176
rect 77260 34628 77300 35848
rect 77356 34712 77396 36763
rect 77452 36728 77492 37351
rect 77452 36679 77492 36688
rect 77547 36140 77589 36149
rect 77547 36100 77548 36140
rect 77588 36100 77589 36140
rect 77547 36091 77589 36100
rect 77548 36006 77588 36091
rect 77452 35888 77492 35897
rect 77452 35645 77492 35848
rect 77644 35888 77684 37948
rect 78508 37568 78548 37577
rect 78124 37400 78164 37409
rect 77931 37232 77973 37241
rect 77931 37192 77932 37232
rect 77972 37192 77973 37232
rect 77931 37183 77973 37192
rect 77932 37098 77972 37183
rect 77644 35839 77684 35848
rect 77836 36056 77876 36065
rect 77451 35636 77493 35645
rect 77451 35596 77452 35636
rect 77492 35596 77493 35636
rect 77451 35587 77493 35596
rect 77643 35384 77685 35393
rect 77643 35344 77644 35384
rect 77684 35344 77685 35384
rect 77643 35335 77685 35344
rect 77451 35216 77493 35225
rect 77451 35176 77452 35216
rect 77492 35176 77493 35216
rect 77451 35167 77493 35176
rect 77452 35082 77492 35167
rect 77356 34672 77588 34712
rect 77260 34579 77300 34588
rect 77452 34544 77492 34553
rect 77356 34504 77452 34544
rect 77356 34460 77396 34504
rect 77452 34495 77492 34504
rect 77164 34420 77396 34460
rect 76972 34327 77012 34336
rect 77452 34376 77492 34385
rect 77548 34376 77588 34672
rect 77644 34385 77684 35335
rect 77836 35225 77876 36016
rect 78124 35477 78164 37360
rect 78316 37400 78356 37411
rect 78508 37409 78548 37528
rect 78316 37325 78356 37360
rect 78507 37400 78549 37409
rect 78507 37360 78508 37400
rect 78548 37360 78549 37400
rect 78507 37351 78549 37360
rect 78220 37316 78260 37325
rect 78220 36737 78260 37276
rect 78315 37316 78357 37325
rect 78315 37276 78316 37316
rect 78356 37276 78357 37316
rect 78315 37267 78357 37276
rect 79467 37316 79509 37325
rect 79467 37276 79468 37316
rect 79508 37276 79509 37316
rect 79467 37267 79509 37276
rect 79468 36896 79508 37267
rect 79468 36847 79508 36856
rect 78219 36728 78261 36737
rect 78219 36688 78220 36728
rect 78260 36688 78261 36728
rect 78219 36679 78261 36688
rect 78316 36728 78356 36737
rect 78316 36065 78356 36688
rect 78315 36056 78357 36065
rect 78315 36016 78316 36056
rect 78356 36016 78357 36056
rect 78315 36007 78357 36016
rect 78123 35468 78165 35477
rect 78123 35428 78124 35468
rect 78164 35428 78165 35468
rect 78123 35419 78165 35428
rect 77835 35216 77877 35225
rect 77835 35176 77836 35216
rect 77876 35176 77877 35216
rect 77835 35167 77877 35176
rect 78124 34637 78164 35419
rect 78316 35216 78356 36007
rect 78316 35167 78356 35176
rect 79468 34964 79508 34973
rect 78123 34628 78165 34637
rect 78123 34588 78124 34628
rect 78164 34588 78165 34628
rect 78123 34579 78165 34588
rect 78028 34544 78068 34553
rect 77740 34504 78028 34544
rect 77492 34336 77588 34376
rect 77643 34376 77685 34385
rect 77643 34336 77644 34376
rect 77684 34336 77685 34376
rect 77452 34327 77492 34336
rect 77643 34327 77685 34336
rect 77740 34376 77780 34504
rect 78028 34495 78068 34504
rect 79468 34385 79508 34924
rect 77740 34327 77780 34336
rect 77931 34376 77973 34385
rect 77931 34336 77932 34376
rect 77972 34336 77973 34376
rect 77931 34327 77973 34336
rect 78123 34376 78165 34385
rect 78123 34336 78124 34376
rect 78164 34336 78165 34376
rect 78123 34327 78165 34336
rect 79467 34376 79509 34385
rect 79467 34336 79468 34376
rect 79508 34336 79509 34376
rect 79467 34327 79509 34336
rect 76875 34292 76917 34301
rect 76875 34252 76876 34292
rect 76916 34252 76917 34292
rect 76875 34243 76917 34252
rect 77355 34292 77397 34301
rect 77355 34252 77356 34292
rect 77396 34252 77397 34292
rect 77355 34243 77397 34252
rect 76492 34168 76820 34208
rect 76352 34040 76720 34049
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 76780 33872 76820 34168
rect 76780 33823 76820 33832
rect 77259 33872 77301 33881
rect 77259 33832 77260 33872
rect 77300 33832 77301 33872
rect 77259 33823 77301 33832
rect 76875 33788 76917 33797
rect 76875 33748 76876 33788
rect 76916 33748 76917 33788
rect 76875 33739 76917 33748
rect 76012 33704 76052 33713
rect 76204 33704 76244 33713
rect 76052 33664 76204 33704
rect 76012 33655 76052 33664
rect 76204 33655 76244 33664
rect 76299 33704 76341 33713
rect 76299 33664 76300 33704
rect 76340 33664 76341 33704
rect 76299 33655 76341 33664
rect 76396 33704 76436 33713
rect 76300 33570 76340 33655
rect 76396 33545 76436 33664
rect 76491 33704 76533 33713
rect 76684 33704 76724 33713
rect 76491 33664 76492 33704
rect 76532 33664 76533 33704
rect 76491 33655 76533 33664
rect 76588 33664 76684 33704
rect 76492 33570 76532 33655
rect 76395 33536 76437 33545
rect 76395 33496 76396 33536
rect 76436 33496 76437 33536
rect 76395 33487 76437 33496
rect 76011 33452 76053 33461
rect 76011 33412 76012 33452
rect 76052 33412 76053 33452
rect 76011 33403 76053 33412
rect 76012 33318 76052 33403
rect 76012 32864 76052 32873
rect 76052 32824 76244 32864
rect 76012 32815 76052 32824
rect 75916 32488 76052 32528
rect 76012 32369 76052 32488
rect 75916 32360 75956 32369
rect 75724 32320 75916 32360
rect 75916 32311 75956 32320
rect 76011 32360 76053 32369
rect 76011 32320 76012 32360
rect 76052 32320 76053 32360
rect 76011 32311 76053 32320
rect 75819 32192 75861 32201
rect 76011 32192 76053 32201
rect 75819 32152 75820 32192
rect 75860 32152 75956 32192
rect 75819 32143 75861 32152
rect 75820 32058 75860 32143
rect 75628 30808 75860 30848
rect 75435 30799 75477 30808
rect 75339 30764 75381 30773
rect 75339 30724 75340 30764
rect 75380 30724 75381 30764
rect 75339 30715 75381 30724
rect 75052 30428 75092 30640
rect 75147 30680 75189 30689
rect 75147 30640 75148 30680
rect 75188 30640 75189 30680
rect 75147 30631 75189 30640
rect 75340 30680 75380 30715
rect 75436 30714 75476 30799
rect 75148 30546 75188 30631
rect 75340 30629 75380 30640
rect 75532 30680 75572 30691
rect 75532 30605 75572 30640
rect 75628 30680 75668 30689
rect 75531 30596 75573 30605
rect 75531 30556 75532 30596
rect 75572 30556 75573 30596
rect 75531 30547 75573 30556
rect 75052 30388 75572 30428
rect 75112 30260 75480 30269
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75112 30211 75480 30220
rect 75435 30092 75477 30101
rect 75532 30092 75572 30388
rect 74956 30052 75380 30092
rect 75051 29924 75093 29933
rect 75051 29884 75052 29924
rect 75092 29884 75093 29924
rect 75051 29875 75093 29884
rect 75052 29790 75092 29875
rect 75340 29840 75380 30052
rect 75435 30052 75436 30092
rect 75476 30052 75572 30092
rect 75628 30092 75668 30640
rect 75820 30101 75860 30808
rect 75724 30092 75764 30101
rect 75628 30052 75724 30092
rect 75435 30043 75477 30052
rect 75724 30043 75764 30052
rect 75819 30092 75861 30101
rect 75819 30052 75820 30092
rect 75860 30052 75861 30092
rect 75819 30043 75861 30052
rect 75340 29791 75380 29800
rect 75436 29840 75476 30043
rect 75627 29924 75669 29933
rect 75916 29924 75956 32152
rect 76011 32152 76012 32192
rect 76052 32152 76053 32192
rect 76011 32143 76053 32152
rect 76108 32192 76148 32201
rect 76012 32058 76052 32143
rect 76012 31604 76052 31613
rect 76108 31604 76148 32152
rect 76204 31697 76244 32824
rect 76588 32705 76628 33664
rect 76684 33655 76724 33664
rect 76876 33704 76916 33739
rect 76876 33653 76916 33664
rect 76971 33704 77013 33713
rect 77260 33704 77300 33823
rect 76971 33664 76972 33704
rect 77012 33664 77204 33704
rect 76971 33655 77013 33664
rect 76972 33570 77012 33655
rect 76779 33452 76821 33461
rect 76779 33412 76780 33452
rect 76820 33412 76821 33452
rect 76779 33403 76821 33412
rect 76587 32696 76629 32705
rect 76587 32656 76588 32696
rect 76628 32656 76629 32696
rect 76587 32647 76629 32656
rect 76352 32528 76720 32537
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76352 32479 76720 32488
rect 76299 32360 76341 32369
rect 76299 32320 76300 32360
rect 76340 32320 76341 32360
rect 76299 32311 76341 32320
rect 76491 32360 76533 32369
rect 76491 32320 76492 32360
rect 76532 32320 76533 32360
rect 76491 32311 76533 32320
rect 76203 31688 76245 31697
rect 76203 31648 76204 31688
rect 76244 31648 76245 31688
rect 76203 31639 76245 31648
rect 76052 31564 76148 31604
rect 76012 31555 76052 31564
rect 76203 31520 76245 31529
rect 76203 31480 76204 31520
rect 76244 31480 76245 31520
rect 76203 31471 76245 31480
rect 76012 31184 76052 31193
rect 76012 30689 76052 31144
rect 76107 31184 76149 31193
rect 76107 31144 76108 31184
rect 76148 31144 76149 31184
rect 76204 31184 76244 31471
rect 76300 31193 76340 32311
rect 76492 31529 76532 32311
rect 76683 32276 76725 32285
rect 76683 32236 76684 32276
rect 76724 32236 76725 32276
rect 76683 32227 76725 32236
rect 76780 32276 76820 33403
rect 77164 33116 77204 33664
rect 77260 33655 77300 33664
rect 77164 32873 77204 33076
rect 77260 33452 77300 33461
rect 77163 32864 77205 32873
rect 77163 32824 77164 32864
rect 77204 32824 77205 32864
rect 77163 32815 77205 32824
rect 76780 32227 76820 32236
rect 77068 32276 77108 32285
rect 77260 32276 77300 33412
rect 77108 32236 77300 32276
rect 77068 32227 77108 32236
rect 76684 32192 76724 32227
rect 76684 32141 76724 32152
rect 76875 32192 76917 32201
rect 76875 32152 76876 32192
rect 76916 32152 76917 32192
rect 76875 32143 76917 32152
rect 76876 32058 76916 32143
rect 76491 31520 76533 31529
rect 76491 31480 76492 31520
rect 76532 31480 76533 31520
rect 77356 31520 77396 34243
rect 77644 34242 77684 34327
rect 77932 34242 77972 34327
rect 78124 34242 78164 34327
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77451 33655 77493 33664
rect 77548 33704 77588 33713
rect 77452 33570 77492 33655
rect 77548 33461 77588 33664
rect 78411 33704 78453 33713
rect 78411 33664 78412 33704
rect 78452 33664 78453 33704
rect 78411 33655 78453 33664
rect 77836 33536 77876 33545
rect 77547 33452 77589 33461
rect 77547 33412 77548 33452
rect 77588 33412 77589 33452
rect 77547 33403 77589 33412
rect 77836 33140 77876 33496
rect 77548 33100 77876 33140
rect 77452 32864 77492 32873
rect 77452 32369 77492 32824
rect 77451 32360 77493 32369
rect 77451 32320 77452 32360
rect 77492 32320 77493 32360
rect 77451 32311 77493 32320
rect 77452 32192 77492 32201
rect 77548 32192 77588 33100
rect 78124 33032 78164 33041
rect 78124 32873 78164 32992
rect 78412 33032 78452 33655
rect 78412 32983 78452 32992
rect 77740 32864 77780 32873
rect 77740 32201 77780 32824
rect 77835 32864 77877 32873
rect 77835 32824 77836 32864
rect 77876 32824 77877 32864
rect 77835 32815 77877 32824
rect 78123 32864 78165 32873
rect 78123 32824 78124 32864
rect 78164 32824 78165 32864
rect 78123 32815 78165 32824
rect 78316 32864 78356 32873
rect 77836 32730 77876 32815
rect 78316 32612 78356 32824
rect 78507 32864 78549 32873
rect 78507 32824 78508 32864
rect 78548 32824 78549 32864
rect 78507 32815 78549 32824
rect 78508 32730 78548 32815
rect 78220 32572 78356 32612
rect 77492 32152 77588 32192
rect 77739 32192 77781 32201
rect 77739 32152 77740 32192
rect 77780 32152 77781 32192
rect 77452 32143 77492 32152
rect 77739 32143 77781 32152
rect 77836 31520 77876 31529
rect 77356 31480 77780 31520
rect 76491 31471 76533 31480
rect 76779 31352 76821 31361
rect 76779 31312 76780 31352
rect 76820 31312 76821 31352
rect 76779 31303 76821 31312
rect 76972 31352 77012 31361
rect 76299 31184 76341 31193
rect 76204 31144 76252 31184
rect 76107 31135 76149 31144
rect 76011 30680 76053 30689
rect 76011 30640 76012 30680
rect 76052 30640 76053 30680
rect 76011 30631 76053 30640
rect 76108 30269 76148 31135
rect 76212 31100 76252 31144
rect 76299 31144 76300 31184
rect 76340 31144 76341 31184
rect 76299 31135 76341 31144
rect 76204 31060 76252 31100
rect 76204 30680 76244 31060
rect 76352 31016 76720 31025
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76352 30967 76720 30976
rect 76491 30764 76533 30773
rect 76491 30724 76492 30764
rect 76532 30724 76533 30764
rect 76491 30715 76533 30724
rect 76107 30260 76149 30269
rect 76107 30220 76108 30260
rect 76148 30220 76149 30260
rect 76107 30211 76149 30220
rect 75627 29884 75628 29924
rect 75668 29884 75669 29924
rect 75627 29875 75669 29884
rect 75724 29884 75956 29924
rect 75436 29791 75476 29800
rect 75531 29840 75573 29849
rect 75531 29800 75532 29840
rect 75572 29800 75573 29840
rect 75531 29791 75573 29800
rect 75532 29706 75572 29791
rect 74859 29672 74901 29681
rect 75244 29672 75284 29681
rect 74859 29632 74860 29672
rect 74900 29632 74901 29672
rect 74859 29623 74901 29632
rect 74956 29632 75244 29672
rect 74860 29538 74900 29623
rect 74668 29119 74708 29128
rect 74956 28580 74996 29632
rect 75244 29623 75284 29632
rect 75112 28748 75480 28757
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75112 28699 75480 28708
rect 75339 28580 75381 28589
rect 74956 28540 75284 28580
rect 75244 28328 75284 28540
rect 75339 28540 75340 28580
rect 75380 28540 75381 28580
rect 75339 28531 75381 28540
rect 75244 28279 75284 28288
rect 75340 28244 75380 28531
rect 75435 28328 75477 28337
rect 75435 28288 75436 28328
rect 75476 28288 75477 28328
rect 75435 28279 75477 28288
rect 75532 28328 75572 28337
rect 75340 28195 75380 28204
rect 75436 28194 75476 28279
rect 75532 27908 75572 28288
rect 75340 27868 75572 27908
rect 75243 27740 75285 27749
rect 75243 27700 75244 27740
rect 75284 27700 75285 27740
rect 75243 27691 75285 27700
rect 74860 27656 74900 27665
rect 74764 27616 74860 27656
rect 74764 26825 74804 27616
rect 74860 27607 74900 27616
rect 75051 27656 75093 27665
rect 75051 27616 75052 27656
rect 75092 27616 75093 27656
rect 75051 27607 75093 27616
rect 75148 27656 75188 27665
rect 75052 27522 75092 27607
rect 74860 27404 74900 27413
rect 75148 27404 75188 27616
rect 75244 27413 75284 27691
rect 74860 26909 74900 27364
rect 74956 27364 75188 27404
rect 75243 27404 75285 27413
rect 75243 27364 75244 27404
rect 75284 27364 75285 27404
rect 75340 27404 75380 27868
rect 75628 27824 75668 29875
rect 75724 29840 75764 29884
rect 76011 29840 76053 29849
rect 75724 29791 75764 29800
rect 75916 29798 75956 29807
rect 75819 29756 75861 29765
rect 75819 29716 75820 29756
rect 75860 29716 75861 29756
rect 75819 29707 75861 29716
rect 76011 29800 76012 29840
rect 76052 29800 76053 29840
rect 76011 29791 76053 29800
rect 75820 29336 75860 29707
rect 75916 29681 75956 29758
rect 76012 29706 76052 29791
rect 75915 29672 75957 29681
rect 75915 29632 75916 29672
rect 75956 29632 75957 29672
rect 75915 29623 75957 29632
rect 75820 29261 75860 29296
rect 75819 29252 75861 29261
rect 75819 29212 75820 29252
rect 75860 29212 75861 29252
rect 75819 29203 75861 29212
rect 75820 29172 75860 29203
rect 76108 29168 76148 29177
rect 76204 29168 76244 30640
rect 76492 30680 76532 30715
rect 76492 30629 76532 30640
rect 76587 30680 76629 30689
rect 76587 30640 76588 30680
rect 76628 30640 76629 30680
rect 76587 30631 76629 30640
rect 76588 30546 76628 30631
rect 76780 30521 76820 31303
rect 76491 30512 76533 30521
rect 76491 30472 76492 30512
rect 76532 30472 76533 30512
rect 76491 30463 76533 30472
rect 76779 30512 76821 30521
rect 76779 30472 76780 30512
rect 76820 30472 76821 30512
rect 76779 30463 76821 30472
rect 76876 30512 76916 30521
rect 76972 30512 77012 31312
rect 77163 31352 77205 31361
rect 77163 31312 77164 31352
rect 77204 31312 77205 31352
rect 77163 31303 77205 31312
rect 77452 31352 77492 31361
rect 77067 31268 77109 31277
rect 77067 31228 77068 31268
rect 77108 31228 77109 31268
rect 77067 31219 77109 31228
rect 77068 31134 77108 31219
rect 77164 31218 77204 31303
rect 77452 31193 77492 31312
rect 77644 31352 77684 31361
rect 77548 31268 77588 31277
rect 77451 31184 77493 31193
rect 77451 31144 77452 31184
rect 77492 31144 77493 31184
rect 77451 31135 77493 31144
rect 77163 31100 77205 31109
rect 77163 31060 77164 31100
rect 77204 31060 77205 31100
rect 77163 31051 77205 31060
rect 76916 30472 77012 30512
rect 77068 30680 77108 30689
rect 76876 30463 76916 30472
rect 76492 29840 76532 30463
rect 77068 30092 77108 30640
rect 77068 30043 77108 30052
rect 76588 30008 76628 30017
rect 76628 29968 76916 30008
rect 76588 29959 76628 29968
rect 76492 29791 76532 29800
rect 76684 29840 76724 29849
rect 76724 29800 76820 29840
rect 76684 29791 76724 29800
rect 76352 29504 76720 29513
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76352 29455 76720 29464
rect 76683 29336 76725 29345
rect 76683 29296 76684 29336
rect 76724 29296 76725 29336
rect 76683 29287 76725 29296
rect 76491 29252 76533 29261
rect 76491 29212 76492 29252
rect 76532 29212 76533 29252
rect 76491 29203 76533 29212
rect 76148 29128 76244 29168
rect 76396 29168 76436 29177
rect 76108 29009 76148 29128
rect 76107 29000 76149 29009
rect 76107 28960 76108 29000
rect 76148 28960 76149 29000
rect 76107 28951 76149 28960
rect 76396 28421 76436 29128
rect 76492 29118 76532 29203
rect 76395 28412 76437 28421
rect 76395 28372 76396 28412
rect 76436 28372 76437 28412
rect 76395 28363 76437 28372
rect 76684 28328 76724 29287
rect 76780 29000 76820 29800
rect 76780 28951 76820 28960
rect 76779 28664 76821 28673
rect 76779 28624 76780 28664
rect 76820 28624 76821 28664
rect 76779 28615 76821 28624
rect 76780 28580 76820 28615
rect 76780 28529 76820 28540
rect 76876 28337 76916 29968
rect 77068 29840 77108 29849
rect 77068 29345 77108 29800
rect 77164 29672 77204 31051
rect 77452 30689 77492 30774
rect 77451 30680 77493 30689
rect 77451 30640 77452 30680
rect 77492 30640 77493 30680
rect 77451 30631 77493 30640
rect 77548 30512 77588 31228
rect 77644 30773 77684 31312
rect 77643 30764 77685 30773
rect 77643 30724 77644 30764
rect 77684 30724 77685 30764
rect 77643 30715 77685 30724
rect 77644 30521 77684 30715
rect 77356 30472 77588 30512
rect 77643 30512 77685 30521
rect 77643 30472 77644 30512
rect 77684 30472 77685 30512
rect 77259 30260 77301 30269
rect 77259 30220 77260 30260
rect 77300 30220 77301 30260
rect 77259 30211 77301 30220
rect 77260 29840 77300 30211
rect 77260 29791 77300 29800
rect 77356 29840 77396 30472
rect 77643 30463 77685 30472
rect 77548 30008 77588 30017
rect 77356 29791 77396 29800
rect 77452 29968 77548 30008
rect 77259 29672 77301 29681
rect 77164 29632 77260 29672
rect 77300 29632 77301 29672
rect 77259 29623 77301 29632
rect 77067 29336 77109 29345
rect 77067 29296 77068 29336
rect 77108 29296 77109 29336
rect 77067 29287 77109 29296
rect 77068 29168 77108 29177
rect 77068 28673 77108 29128
rect 77067 28664 77109 28673
rect 77067 28624 77068 28664
rect 77108 28624 77109 28664
rect 77067 28615 77109 28624
rect 76780 28328 76820 28337
rect 76684 28288 76780 28328
rect 76780 28279 76820 28288
rect 76875 28328 76917 28337
rect 76972 28328 77012 28337
rect 76875 28288 76876 28328
rect 76916 28288 76972 28328
rect 76875 28279 76917 28288
rect 76972 28279 77012 28288
rect 77068 28328 77108 28337
rect 76876 28194 76916 28279
rect 77068 28160 77108 28288
rect 77260 28328 77300 29623
rect 77452 29168 77492 29968
rect 77548 29959 77588 29968
rect 77452 29119 77492 29128
rect 77260 28279 77300 28288
rect 77451 28328 77493 28337
rect 77451 28288 77452 28328
rect 77492 28288 77493 28328
rect 77451 28279 77493 28288
rect 77356 28244 77396 28253
rect 77356 28160 77396 28204
rect 77452 28194 77492 28279
rect 77068 28120 77396 28160
rect 76352 27992 76720 28001
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76352 27943 76720 27952
rect 75532 27784 75668 27824
rect 75435 27740 75477 27749
rect 75435 27700 75436 27740
rect 75476 27700 75477 27740
rect 75435 27691 75477 27700
rect 75436 27656 75476 27691
rect 75436 27605 75476 27616
rect 75436 27404 75476 27413
rect 75340 27364 75436 27404
rect 74859 26900 74901 26909
rect 74859 26860 74860 26900
rect 74900 26860 74901 26900
rect 74859 26851 74901 26860
rect 74763 26816 74805 26825
rect 74763 26776 74764 26816
rect 74804 26776 74805 26816
rect 74763 26767 74805 26776
rect 74763 26396 74805 26405
rect 74763 26356 74764 26396
rect 74804 26356 74805 26396
rect 74763 26347 74805 26356
rect 74667 26312 74709 26321
rect 74667 26272 74668 26312
rect 74708 26272 74709 26312
rect 74667 26263 74709 26272
rect 74668 26178 74708 26263
rect 74764 26144 74804 26347
rect 74956 26312 74996 27364
rect 75243 27355 75285 27364
rect 75436 27355 75476 27364
rect 75112 27236 75480 27245
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75112 27187 75480 27196
rect 75147 27068 75189 27077
rect 75147 27028 75148 27068
rect 75188 27028 75189 27068
rect 75147 27019 75189 27028
rect 75339 27068 75381 27077
rect 75339 27028 75340 27068
rect 75380 27028 75381 27068
rect 75339 27019 75381 27028
rect 74956 26272 75092 26312
rect 74859 26228 74901 26237
rect 74859 26188 74860 26228
rect 74900 26188 74901 26228
rect 74859 26179 74901 26188
rect 74764 26095 74804 26104
rect 74860 26144 74900 26179
rect 74860 26093 74900 26104
rect 74956 26144 74996 26153
rect 74859 25976 74901 25985
rect 74956 25976 74996 26104
rect 74859 25936 74860 25976
rect 74900 25936 74996 25976
rect 75052 25976 75092 26272
rect 75148 26144 75188 27019
rect 75148 26095 75188 26104
rect 75244 26228 75284 26237
rect 75244 25976 75284 26188
rect 75052 25936 75284 25976
rect 75340 26144 75380 27019
rect 75435 26900 75477 26909
rect 75435 26860 75436 26900
rect 75476 26860 75477 26900
rect 75435 26851 75477 26860
rect 75436 26766 75476 26851
rect 74859 25927 74901 25936
rect 75340 25892 75380 26104
rect 75436 26144 75476 26153
rect 75436 25985 75476 26104
rect 75435 25976 75477 25985
rect 75435 25936 75436 25976
rect 75476 25936 75477 25976
rect 75435 25927 75477 25936
rect 74956 25852 75380 25892
rect 74572 25348 74708 25388
rect 74475 25304 74517 25313
rect 74380 25264 74476 25304
rect 74516 25264 74517 25304
rect 74475 25255 74517 25264
rect 74476 25170 74516 25255
rect 74571 25220 74613 25229
rect 74571 25180 74572 25220
rect 74612 25180 74613 25220
rect 74571 25171 74613 25180
rect 74380 24800 74420 24809
rect 74188 24760 74380 24800
rect 74380 24751 74420 24760
rect 74475 24800 74517 24809
rect 74475 24760 74476 24800
rect 74516 24760 74517 24800
rect 74475 24751 74517 24760
rect 74284 24632 74324 24641
rect 74092 24592 74284 24632
rect 74284 24583 74324 24592
rect 74476 24632 74516 24751
rect 74476 24583 74516 24592
rect 74572 24632 74612 25171
rect 74572 24583 74612 24592
rect 74668 24464 74708 25348
rect 74956 24809 74996 25852
rect 75112 25724 75480 25733
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75112 25675 75480 25684
rect 75435 25388 75477 25397
rect 75435 25348 75436 25388
rect 75476 25348 75477 25388
rect 75435 25339 75477 25348
rect 74955 24800 74997 24809
rect 74955 24760 74956 24800
rect 74996 24760 74997 24800
rect 74955 24751 74997 24760
rect 75436 24632 75476 25339
rect 75436 24583 75476 24592
rect 74092 24424 74708 24464
rect 73803 23960 73845 23969
rect 73803 23920 73804 23960
rect 73844 23920 73845 23960
rect 73803 23911 73845 23920
rect 73995 23960 74037 23969
rect 73995 23920 73996 23960
rect 74036 23920 74037 23960
rect 73995 23911 74037 23920
rect 74092 23792 74132 24424
rect 73748 23752 74036 23792
rect 73708 23743 73748 23752
rect 73804 23624 73844 23633
rect 73804 23060 73844 23584
rect 73996 23060 74036 23752
rect 74092 23743 74132 23752
rect 74188 23624 74228 23633
rect 74188 23060 74228 23584
rect 74380 23060 74420 24424
rect 75243 24212 75285 24221
rect 75243 24172 75244 24212
rect 75284 24172 75285 24212
rect 75243 24163 75285 24172
rect 74475 24044 74517 24053
rect 74475 24004 74476 24044
rect 74516 24004 74517 24044
rect 74475 23995 74517 24004
rect 74476 23792 74516 23995
rect 74859 23960 74901 23969
rect 74859 23920 74860 23960
rect 74900 23920 74901 23960
rect 74859 23911 74901 23920
rect 74476 23297 74516 23752
rect 74860 23792 74900 23911
rect 74572 23624 74612 23633
rect 74475 23288 74517 23297
rect 74475 23248 74476 23288
rect 74516 23248 74517 23288
rect 74475 23239 74517 23248
rect 74572 23060 74612 23584
rect 74860 23465 74900 23752
rect 75244 23792 75284 24163
rect 75532 23792 75572 27784
rect 75628 27656 75668 27665
rect 75628 27077 75668 27616
rect 75724 27656 75764 27665
rect 75627 27068 75669 27077
rect 75627 27028 75628 27068
rect 75668 27028 75669 27068
rect 75627 27019 75669 27028
rect 75724 26993 75764 27616
rect 76684 27656 76724 27665
rect 75723 26984 75765 26993
rect 75723 26944 75724 26984
rect 75764 26944 75765 26984
rect 75723 26935 75765 26944
rect 75627 26816 75669 26825
rect 75627 26776 75628 26816
rect 75668 26776 75669 26816
rect 75627 26767 75669 26776
rect 75724 26816 75764 26825
rect 75628 26682 75668 26767
rect 75627 26564 75669 26573
rect 75627 26524 75628 26564
rect 75668 26524 75669 26564
rect 75627 26515 75669 26524
rect 75628 26228 75668 26515
rect 75724 26405 75764 26776
rect 75820 26816 75860 26825
rect 75723 26396 75765 26405
rect 75723 26356 75724 26396
rect 75764 26356 75765 26396
rect 75723 26347 75765 26356
rect 75820 26237 75860 26776
rect 75915 26816 75957 26825
rect 75915 26776 75916 26816
rect 75956 26776 75957 26816
rect 75915 26767 75957 26776
rect 76204 26816 76244 26825
rect 75916 26682 75956 26767
rect 76204 26657 76244 26776
rect 76492 26816 76532 26825
rect 76492 26657 76532 26776
rect 76587 26816 76629 26825
rect 76587 26776 76588 26816
rect 76628 26776 76629 26816
rect 76587 26767 76629 26776
rect 76588 26682 76628 26767
rect 76203 26648 76245 26657
rect 76203 26608 76204 26648
rect 76244 26608 76245 26648
rect 76203 26599 76245 26608
rect 76491 26648 76533 26657
rect 76491 26608 76492 26648
rect 76532 26608 76533 26648
rect 76684 26648 76724 27616
rect 76779 27656 76821 27665
rect 76779 27616 76780 27656
rect 76820 27616 76821 27656
rect 76779 27607 76821 27616
rect 76876 27656 76916 27665
rect 76780 27522 76820 27607
rect 76876 27068 76916 27616
rect 76971 27656 77013 27665
rect 76971 27616 76972 27656
rect 77012 27616 77013 27656
rect 76971 27607 77013 27616
rect 77164 27656 77204 27665
rect 76876 27019 76916 27028
rect 76684 26608 76820 26648
rect 76491 26599 76533 26608
rect 76352 26480 76720 26489
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76352 26431 76720 26440
rect 76780 26312 76820 26608
rect 76684 26272 76820 26312
rect 76875 26312 76917 26321
rect 76875 26272 76876 26312
rect 76916 26272 76917 26312
rect 75819 26228 75861 26237
rect 75628 26188 75764 26228
rect 75627 25976 75669 25985
rect 75627 25936 75628 25976
rect 75668 25936 75669 25976
rect 75627 25927 75669 25936
rect 75628 25556 75668 25927
rect 75628 25507 75668 25516
rect 75724 25397 75764 26188
rect 75819 26188 75820 26228
rect 75860 26188 75861 26228
rect 75819 26179 75861 26188
rect 75915 26144 75957 26153
rect 75915 26104 75916 26144
rect 75956 26104 75957 26144
rect 75915 26095 75957 26104
rect 76395 26144 76437 26153
rect 76395 26104 76396 26144
rect 76436 26104 76437 26144
rect 76395 26095 76437 26104
rect 75819 25976 75861 25985
rect 75819 25936 75820 25976
rect 75860 25936 75861 25976
rect 75819 25927 75861 25936
rect 75723 25388 75765 25397
rect 75723 25348 75724 25388
rect 75764 25348 75765 25388
rect 75723 25339 75765 25348
rect 75820 25304 75860 25927
rect 75916 25472 75956 26095
rect 76203 25892 76245 25901
rect 76203 25852 76204 25892
rect 76244 25852 76245 25892
rect 76203 25843 76245 25852
rect 75916 25423 75956 25432
rect 75820 25255 75860 25264
rect 76012 25305 76052 25313
rect 76012 25304 76148 25305
rect 76052 25265 76148 25304
rect 76052 25264 76053 25265
rect 76012 25255 76052 25264
rect 75628 25136 75668 25145
rect 75668 25096 75860 25136
rect 75628 25087 75668 25096
rect 75820 24716 75860 25096
rect 75820 24667 75860 24676
rect 75723 24632 75765 24641
rect 75723 24592 75724 24632
rect 75764 24592 75765 24632
rect 75723 24583 75765 24592
rect 75724 24498 75764 24583
rect 76108 24464 76148 25265
rect 76204 25304 76244 25843
rect 76204 24977 76244 25264
rect 76300 25229 76340 25314
rect 76396 25304 76436 26095
rect 76684 25985 76724 26272
rect 76875 26263 76917 26272
rect 76876 26178 76916 26263
rect 76780 26144 76820 26153
rect 76683 25976 76725 25985
rect 76683 25936 76684 25976
rect 76724 25936 76725 25976
rect 76683 25927 76725 25936
rect 76780 25901 76820 26104
rect 76972 26144 77012 27607
rect 77164 27497 77204 27616
rect 77356 27656 77396 27665
rect 77163 27488 77205 27497
rect 77163 27448 77164 27488
rect 77204 27448 77205 27488
rect 77163 27439 77205 27448
rect 77260 27404 77300 27413
rect 77068 26732 77108 26741
rect 77068 26321 77108 26692
rect 77067 26312 77109 26321
rect 77067 26272 77068 26312
rect 77108 26272 77109 26312
rect 77067 26263 77109 26272
rect 76972 26095 77012 26104
rect 77068 26144 77108 26153
rect 77260 26144 77300 27364
rect 77356 26657 77396 27616
rect 77548 27488 77588 27497
rect 77452 26816 77492 26825
rect 77548 26816 77588 27448
rect 77492 26776 77588 26816
rect 77452 26767 77492 26776
rect 77355 26648 77397 26657
rect 77355 26608 77356 26648
rect 77396 26608 77397 26648
rect 77355 26599 77397 26608
rect 77108 26104 77300 26144
rect 77068 26095 77108 26104
rect 77740 26060 77780 31480
rect 77836 30689 77876 31480
rect 78220 31361 78260 32572
rect 78316 32192 78356 32201
rect 78316 31697 78356 32152
rect 79467 32192 79509 32201
rect 79467 32152 79468 32192
rect 79508 32152 79509 32192
rect 79467 32143 79509 32152
rect 79468 32108 79508 32143
rect 79468 32057 79508 32068
rect 78315 31688 78357 31697
rect 78315 31648 78316 31688
rect 78356 31648 78357 31688
rect 78315 31639 78357 31648
rect 78219 31352 78261 31361
rect 78219 31312 78220 31352
rect 78260 31312 78261 31352
rect 78219 31303 78261 31312
rect 77835 30680 77877 30689
rect 77835 30640 77836 30680
rect 77876 30640 77877 30680
rect 77835 30631 77877 30640
rect 78316 30680 78356 31639
rect 77835 30512 77877 30521
rect 77835 30472 77836 30512
rect 77876 30472 77877 30512
rect 77835 30463 77877 30472
rect 77836 28757 77876 30463
rect 78316 29168 78356 30640
rect 79467 30512 79509 30521
rect 79467 30472 79468 30512
rect 79508 30472 79509 30512
rect 79467 30463 79509 30472
rect 79468 30378 79508 30463
rect 78316 29119 78356 29128
rect 79468 28916 79508 28925
rect 77835 28748 77877 28757
rect 77835 28708 77836 28748
rect 77876 28708 77877 28748
rect 77835 28699 77877 28708
rect 79468 28337 79508 28876
rect 78123 28328 78165 28337
rect 78123 28288 78124 28328
rect 78164 28288 78165 28328
rect 78123 28279 78165 28288
rect 79467 28328 79509 28337
rect 79467 28288 79468 28328
rect 79508 28288 79509 28328
rect 79467 28279 79509 28288
rect 77260 26020 77780 26060
rect 76779 25892 76821 25901
rect 76779 25852 76780 25892
rect 76820 25852 76821 25892
rect 76779 25843 76821 25852
rect 76588 25432 76820 25472
rect 76396 25255 76436 25264
rect 76492 25304 76532 25313
rect 76588 25304 76628 25432
rect 76532 25264 76628 25304
rect 76492 25255 76532 25264
rect 76684 25229 76724 25314
rect 76299 25220 76341 25229
rect 76299 25180 76300 25220
rect 76340 25180 76341 25220
rect 76299 25171 76341 25180
rect 76683 25220 76725 25229
rect 76683 25180 76684 25220
rect 76724 25180 76725 25220
rect 76683 25171 76725 25180
rect 76203 24968 76245 24977
rect 76203 24928 76204 24968
rect 76244 24928 76245 24968
rect 76203 24919 76245 24928
rect 76352 24968 76720 24977
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76352 24919 76720 24928
rect 76491 24800 76533 24809
rect 76780 24800 76820 25432
rect 77068 25304 77108 25313
rect 77108 25264 77204 25304
rect 77068 25255 77108 25264
rect 76491 24760 76492 24800
rect 76532 24760 76533 24800
rect 76491 24751 76533 24760
rect 76588 24760 76820 24800
rect 76492 24632 76532 24751
rect 76588 24716 76628 24760
rect 76588 24667 76628 24676
rect 76492 24583 76532 24592
rect 76683 24632 76725 24641
rect 76683 24592 76684 24632
rect 76724 24592 76725 24632
rect 76683 24583 76725 24592
rect 76684 24498 76724 24583
rect 76108 24415 76148 24424
rect 77164 24464 77204 25264
rect 77164 24415 77204 24424
rect 75628 23792 75668 23801
rect 76107 23792 76149 23801
rect 75532 23752 75628 23792
rect 75668 23752 75860 23792
rect 75244 23633 75284 23752
rect 75628 23743 75668 23752
rect 75820 23708 75860 23752
rect 76107 23752 76108 23792
rect 76148 23752 76149 23792
rect 76107 23743 76149 23752
rect 76491 23792 76533 23801
rect 76491 23752 76492 23792
rect 76532 23752 76533 23792
rect 76491 23743 76533 23752
rect 76971 23792 77013 23801
rect 76971 23752 76972 23792
rect 77012 23752 77013 23792
rect 76971 23743 77013 23752
rect 77260 23792 77300 26020
rect 77835 25892 77877 25901
rect 77835 25852 77836 25892
rect 77876 25852 77877 25892
rect 77835 25843 77877 25852
rect 75820 23668 76052 23708
rect 74956 23624 74996 23633
rect 74859 23456 74901 23465
rect 74859 23416 74860 23456
rect 74900 23416 74901 23456
rect 74859 23407 74901 23416
rect 74859 23288 74901 23297
rect 74859 23248 74860 23288
rect 74900 23248 74901 23288
rect 74859 23239 74901 23248
rect 73612 23020 73695 23060
rect 73804 23020 73940 23060
rect 73996 23020 74095 23060
rect 74188 23020 74324 23060
rect 74380 23020 74495 23060
rect 74572 23020 74785 23060
rect 73516 22744 73585 22784
rect 73545 22596 73585 22744
rect 73655 22596 73695 23020
rect 73900 22784 73940 23020
rect 73900 22744 73985 22784
rect 73945 22596 73985 22744
rect 74055 22596 74095 23020
rect 74284 22784 74324 23020
rect 74284 22744 74385 22784
rect 74345 22596 74385 22744
rect 74455 22596 74495 23020
rect 74745 22596 74785 23020
rect 74860 22868 74900 23239
rect 74855 22828 74900 22868
rect 74855 22596 74895 22828
rect 74956 22784 74996 23584
rect 75243 23624 75285 23633
rect 75243 23584 75244 23624
rect 75284 23584 75285 23624
rect 75243 23575 75285 23584
rect 75340 23624 75380 23633
rect 75243 23456 75285 23465
rect 75243 23416 75244 23456
rect 75284 23416 75285 23456
rect 75243 23407 75285 23416
rect 75244 23060 75284 23407
rect 75340 23060 75380 23584
rect 75627 23624 75669 23633
rect 75627 23584 75628 23624
rect 75668 23584 75669 23624
rect 75627 23575 75669 23584
rect 75724 23624 75764 23633
rect 75764 23584 75956 23624
rect 75724 23575 75764 23584
rect 75628 23060 75668 23575
rect 75244 23020 75295 23060
rect 75340 23020 75585 23060
rect 75628 23020 75695 23060
rect 74956 22744 75185 22784
rect 75145 22596 75185 22744
rect 75255 22596 75295 23020
rect 75545 22596 75585 23020
rect 75655 22596 75695 23020
rect 75916 22784 75956 23584
rect 76012 23060 76052 23668
rect 76108 23658 76148 23743
rect 76204 23624 76244 23633
rect 76204 23060 76244 23584
rect 76492 23060 76532 23743
rect 76876 23624 76916 23633
rect 76780 23584 76876 23624
rect 76780 23060 76820 23584
rect 76876 23575 76916 23584
rect 76972 23060 77012 23743
rect 77164 23624 77204 23633
rect 77164 23060 77204 23584
rect 77260 23060 77300 23752
rect 77451 23792 77493 23801
rect 77740 23792 77780 23801
rect 77836 23792 77876 25843
rect 77931 25304 77973 25313
rect 77931 25264 77932 25304
rect 77972 25264 77973 25304
rect 77931 25255 77973 25264
rect 77932 25170 77972 25255
rect 78124 23792 78164 28279
rect 78316 26816 78356 26825
rect 78316 25313 78356 26776
rect 78507 26648 78549 26657
rect 78507 26608 78508 26648
rect 78548 26608 78549 26648
rect 78507 26599 78549 26608
rect 79467 26648 79509 26657
rect 79467 26608 79468 26648
rect 79508 26608 79509 26648
rect 79467 26599 79509 26608
rect 78315 25304 78357 25313
rect 78315 25264 78316 25304
rect 78356 25264 78357 25304
rect 78315 25255 78357 25264
rect 78508 23792 78548 26599
rect 79468 26514 79508 26599
rect 79084 25136 79124 25145
rect 78988 25096 79084 25136
rect 78988 24641 79028 25096
rect 79084 25087 79124 25096
rect 78987 24632 79029 24641
rect 78987 24592 78988 24632
rect 79028 24592 79029 24632
rect 78987 24583 79029 24592
rect 77451 23752 77452 23792
rect 77492 23752 77684 23792
rect 77451 23743 77493 23752
rect 77452 23658 77492 23743
rect 77548 23624 77588 23633
rect 77548 23060 77588 23584
rect 76012 23020 76095 23060
rect 76204 23020 76340 23060
rect 75916 22744 75985 22784
rect 75945 22596 75985 22744
rect 76055 22596 76095 23020
rect 76300 22784 76340 23020
rect 76455 23020 76532 23060
rect 76745 23020 76820 23060
rect 76876 23020 77012 23060
rect 77145 23020 77204 23060
rect 77255 23020 77300 23060
rect 77545 23020 77588 23060
rect 77644 23060 77684 23752
rect 77780 23752 78068 23792
rect 77740 23743 77780 23752
rect 77836 23624 77876 23633
rect 77836 23060 77876 23584
rect 78028 23060 78068 23752
rect 78164 23752 78452 23792
rect 78124 23743 78164 23752
rect 78220 23624 78260 23633
rect 78220 23060 78260 23584
rect 77644 23020 77695 23060
rect 77836 23020 77985 23060
rect 78028 23020 78095 23060
rect 78220 23020 78356 23060
rect 76300 22744 76385 22784
rect 76345 22596 76385 22744
rect 76455 22596 76495 23020
rect 76745 22596 76785 23020
rect 76876 22784 76916 23020
rect 76855 22744 76916 22784
rect 76855 22596 76895 22744
rect 77145 22596 77185 23020
rect 77255 22596 77295 23020
rect 77545 22596 77585 23020
rect 77655 22596 77695 23020
rect 77945 22596 77985 23020
rect 78055 22596 78095 23020
rect 78316 22784 78356 23020
rect 78412 22868 78452 23752
rect 78508 23060 78548 23752
rect 78796 23792 78836 23801
rect 78988 23792 79028 24583
rect 78836 23752 79028 23792
rect 79083 23792 79125 23801
rect 79083 23752 79084 23792
rect 79124 23752 79125 23792
rect 78604 23624 78644 23633
rect 78644 23584 78740 23624
rect 78604 23575 78644 23584
rect 78700 23060 78740 23584
rect 78796 23465 78836 23752
rect 79083 23743 79125 23752
rect 79372 23792 79412 23801
rect 79084 23658 79124 23743
rect 78892 23624 78932 23633
rect 78795 23456 78837 23465
rect 78795 23416 78796 23456
rect 78836 23416 78837 23456
rect 78795 23407 78837 23416
rect 78892 23060 78932 23584
rect 79180 23624 79220 23633
rect 79372 23624 79412 23752
rect 79220 23584 79412 23624
rect 79180 23575 79220 23584
rect 79275 23456 79317 23465
rect 79275 23416 79276 23456
rect 79316 23416 79317 23456
rect 79275 23407 79317 23416
rect 79276 23060 79316 23407
rect 78508 23020 78644 23060
rect 78700 23020 78785 23060
rect 78892 23020 79185 23060
rect 78412 22828 78495 22868
rect 78316 22744 78385 22784
rect 78345 22596 78385 22744
rect 78455 22596 78495 22828
rect 78604 22793 78644 23020
rect 78603 22784 78645 22793
rect 78603 22744 78604 22784
rect 78644 22744 78645 22784
rect 78603 22735 78645 22744
rect 78745 22596 78785 23020
rect 78854 22784 78896 22793
rect 78854 22744 78855 22784
rect 78895 22744 78896 22784
rect 78854 22735 78896 22744
rect 78855 22596 78895 22735
rect 79145 22596 79185 23020
rect 79255 23020 79316 23060
rect 79372 23060 79412 23584
rect 79468 23624 79508 23633
rect 79508 23584 79700 23624
rect 79468 23575 79508 23584
rect 79660 23060 79700 23584
rect 79372 23020 79585 23060
rect 79255 22596 79295 23020
rect 79545 22596 79585 23020
rect 79655 23020 79700 23060
rect 79655 22596 79695 23020
rect 52971 22028 53013 22037
rect 52971 21988 52972 22028
rect 53012 21988 53013 22028
rect 52971 21979 53013 21988
rect 52724 21568 52916 21608
rect 52684 21559 52724 21568
rect 52588 20189 52628 21559
rect 52684 21020 52724 21029
rect 52972 21020 53012 21979
rect 52724 20980 53012 21020
rect 52684 20971 52724 20980
rect 52587 20180 52629 20189
rect 52587 20140 52588 20180
rect 52628 20140 52629 20180
rect 52587 20131 52629 20140
rect 52299 18584 52341 18593
rect 52684 18584 52724 18593
rect 52299 18544 52300 18584
rect 52340 18544 52341 18584
rect 52299 18535 52341 18544
rect 52492 18544 52684 18584
rect 52300 18450 52340 18535
rect 52396 18332 52436 18341
rect 52396 17333 52436 18292
rect 52395 17324 52437 17333
rect 52395 17284 52396 17324
rect 52436 17284 52437 17324
rect 52395 17275 52437 17284
rect 52492 17165 52532 18544
rect 52684 18535 52724 18544
rect 52588 18332 52628 18341
rect 52628 18292 53012 18332
rect 52588 18283 52628 18292
rect 52779 18164 52821 18173
rect 52779 18124 52780 18164
rect 52820 18124 52821 18164
rect 52779 18115 52821 18124
rect 52684 17576 52724 17585
rect 52684 17249 52724 17536
rect 52683 17240 52725 17249
rect 52683 17200 52684 17240
rect 52724 17200 52725 17240
rect 52683 17191 52725 17200
rect 52299 17156 52341 17165
rect 52299 17116 52300 17156
rect 52340 17116 52341 17156
rect 52299 17107 52341 17116
rect 52491 17156 52533 17165
rect 52491 17116 52492 17156
rect 52532 17116 52533 17156
rect 52491 17107 52533 17116
rect 52203 17072 52245 17081
rect 52203 17032 52204 17072
rect 52244 17032 52245 17072
rect 52203 17023 52245 17032
rect 52300 17072 52340 17107
rect 52300 17021 52340 17032
rect 52395 16988 52437 16997
rect 52395 16948 52396 16988
rect 52436 16948 52437 16988
rect 52395 16939 52437 16948
rect 52396 16854 52436 16939
rect 52492 16904 52532 17107
rect 52588 17081 52628 17166
rect 52587 17072 52629 17081
rect 52587 17032 52588 17072
rect 52628 17032 52629 17072
rect 52587 17023 52629 17032
rect 52684 16904 52724 16913
rect 52492 16864 52684 16904
rect 52684 16855 52724 16864
rect 52203 16820 52245 16829
rect 52203 16780 52204 16820
rect 52244 16780 52245 16820
rect 52203 16771 52245 16780
rect 52204 15560 52244 16771
rect 52780 16736 52820 18115
rect 52972 17324 53012 18292
rect 54455 17758 54495 17808
rect 54445 17718 54495 17758
rect 54445 17576 54485 17718
rect 54437 17536 54485 17576
rect 53545 17324 53585 17472
rect 52972 17284 53585 17324
rect 53655 17165 53695 17472
rect 53945 17324 53985 17472
rect 53932 17284 53985 17324
rect 53835 17240 53877 17249
rect 53835 17200 53836 17240
rect 53876 17200 53877 17240
rect 53835 17191 53877 17200
rect 53654 17156 53696 17165
rect 53654 17116 53655 17156
rect 53695 17116 53696 17156
rect 53654 17107 53696 17116
rect 52684 16696 52820 16736
rect 52588 16232 52628 16241
rect 52684 16232 52724 16696
rect 53836 16577 53876 17191
rect 53932 17081 53972 17284
rect 54055 17165 54095 17472
rect 54345 17249 54385 17472
rect 54437 17333 54477 17536
rect 54436 17324 54478 17333
rect 54436 17284 54437 17324
rect 54477 17284 54478 17324
rect 54436 17275 54478 17284
rect 54344 17240 54386 17249
rect 54344 17200 54345 17240
rect 54385 17200 54386 17240
rect 54344 17191 54386 17200
rect 54054 17156 54096 17165
rect 54054 17116 54055 17156
rect 54095 17116 54096 17156
rect 54054 17107 54096 17116
rect 54507 17156 54549 17165
rect 54507 17116 54508 17156
rect 54548 17116 54549 17156
rect 54507 17107 54549 17116
rect 53931 17072 53973 17081
rect 53931 17032 53932 17072
rect 53972 17032 53973 17072
rect 53931 17023 53973 17032
rect 54411 17072 54453 17081
rect 54411 17032 54412 17072
rect 54452 17032 54453 17072
rect 54411 17023 54453 17032
rect 53835 16568 53877 16577
rect 53835 16528 53836 16568
rect 53876 16528 53877 16568
rect 53835 16519 53877 16528
rect 53164 16400 53204 16409
rect 53644 16400 53684 16409
rect 52876 16360 53164 16400
rect 52628 16192 52724 16232
rect 52779 16232 52821 16241
rect 52779 16192 52780 16232
rect 52820 16192 52821 16232
rect 52588 15896 52628 16192
rect 52779 16183 52821 16192
rect 52876 16232 52916 16360
rect 53164 16351 53204 16360
rect 53548 16360 53644 16400
rect 52876 16183 52916 16192
rect 53068 16232 53108 16241
rect 53108 16192 53204 16232
rect 53068 16183 53108 16192
rect 52780 16098 52820 16183
rect 52684 16064 52724 16073
rect 52684 15980 52724 16024
rect 52684 15940 52820 15980
rect 52588 15856 52724 15896
rect 52492 15560 52532 15569
rect 52244 15520 52340 15560
rect 52204 15511 52244 15520
rect 52108 15352 52244 15392
rect 52012 14468 52052 14680
rect 52107 14468 52149 14477
rect 52012 14428 52108 14468
rect 52148 14428 52149 14468
rect 52107 14419 52149 14428
rect 52108 14216 52148 14419
rect 52204 14225 52244 15352
rect 52300 14729 52340 15520
rect 52492 15317 52532 15520
rect 52587 15560 52629 15569
rect 52587 15520 52588 15560
rect 52628 15520 52629 15560
rect 52587 15511 52629 15520
rect 52588 15426 52628 15511
rect 52491 15308 52533 15317
rect 52491 15268 52492 15308
rect 52532 15268 52533 15308
rect 52491 15259 52533 15268
rect 52299 14720 52341 14729
rect 52299 14680 52300 14720
rect 52340 14680 52341 14720
rect 52299 14671 52341 14680
rect 52684 14561 52724 15856
rect 52780 15737 52820 15940
rect 53164 15905 53204 16192
rect 53269 16219 53309 16228
rect 52971 15896 53013 15905
rect 52971 15856 52972 15896
rect 53012 15856 53013 15896
rect 52971 15847 53013 15856
rect 53163 15896 53205 15905
rect 53163 15856 53164 15896
rect 53204 15856 53205 15896
rect 53163 15847 53205 15856
rect 52779 15728 52821 15737
rect 52779 15688 52780 15728
rect 52820 15688 52821 15728
rect 52779 15679 52821 15688
rect 52972 15560 53012 15847
rect 53269 15812 53309 16179
rect 53451 15896 53493 15905
rect 53451 15856 53452 15896
rect 53492 15856 53493 15896
rect 53451 15847 53493 15856
rect 53269 15772 53396 15812
rect 53163 15728 53205 15737
rect 53163 15688 53164 15728
rect 53204 15688 53205 15728
rect 53163 15679 53205 15688
rect 53164 15644 53204 15679
rect 53164 15593 53204 15604
rect 52972 15520 53108 15560
rect 52876 15308 52916 15317
rect 52683 14552 52725 14561
rect 52683 14512 52684 14552
rect 52724 14512 52725 14552
rect 52683 14503 52725 14512
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 52108 14167 52148 14176
rect 52203 14216 52245 14225
rect 52203 14176 52204 14216
rect 52244 14176 52245 14216
rect 52203 14167 52245 14176
rect 52588 14048 52628 14057
rect 52588 12980 52628 14008
rect 52876 14048 52916 15268
rect 52971 14132 53013 14141
rect 52971 14092 52972 14132
rect 53012 14092 53013 14132
rect 52971 14083 53013 14092
rect 52876 13999 52916 14008
rect 52972 13998 53012 14083
rect 53068 14048 53108 15520
rect 53163 15476 53205 15485
rect 53163 15436 53164 15476
rect 53204 15436 53205 15476
rect 53163 15427 53205 15436
rect 53164 14972 53204 15427
rect 53356 15317 53396 15772
rect 53355 15308 53397 15317
rect 53355 15268 53356 15308
rect 53396 15268 53397 15308
rect 53355 15259 53397 15268
rect 53164 14923 53204 14932
rect 53164 14552 53204 14561
rect 53204 14512 53396 14552
rect 53164 14503 53204 14512
rect 53068 13889 53108 14008
rect 53356 14048 53396 14512
rect 53356 13999 53396 14008
rect 53452 14048 53492 15847
rect 53548 15560 53588 16360
rect 53644 16351 53684 16360
rect 54412 16232 54452 17023
rect 54508 16484 54548 17107
rect 54745 17081 54785 17472
rect 54855 17249 54895 17472
rect 55145 17249 55185 17472
rect 54854 17240 54896 17249
rect 54854 17200 54855 17240
rect 54895 17200 54896 17240
rect 54854 17191 54896 17200
rect 55144 17240 55186 17249
rect 55144 17200 55145 17240
rect 55185 17200 55186 17240
rect 55144 17191 55186 17200
rect 54744 17072 54786 17081
rect 55255 17072 55295 17472
rect 55545 17156 55585 17472
rect 54744 17032 54745 17072
rect 54785 17032 54786 17072
rect 54744 17023 54786 17032
rect 54892 17032 55295 17072
rect 55468 17116 55585 17156
rect 54508 16435 54548 16444
rect 54892 16484 54932 17032
rect 55468 16745 55508 17116
rect 55655 17072 55695 17472
rect 55945 17156 55985 17472
rect 55945 17116 55988 17156
rect 55564 17032 55695 17072
rect 55467 16736 55509 16745
rect 55467 16696 55468 16736
rect 55508 16696 55509 16736
rect 55467 16687 55509 16696
rect 54892 16435 54932 16444
rect 55468 16316 55508 16687
rect 55276 16276 55508 16316
rect 54412 16183 54452 16192
rect 54795 16232 54837 16241
rect 54795 16192 54796 16232
rect 54836 16192 54837 16232
rect 54795 16183 54837 16192
rect 55276 16232 55316 16276
rect 55276 16183 55316 16192
rect 54796 16098 54836 16183
rect 55372 16148 55412 16157
rect 55564 16148 55604 17032
rect 55948 16661 55988 17116
rect 56055 17072 56095 17472
rect 56345 17156 56385 17472
rect 56044 17032 56095 17072
rect 56140 17116 56385 17156
rect 55659 16652 55701 16661
rect 55659 16612 55660 16652
rect 55700 16612 55701 16652
rect 55659 16603 55701 16612
rect 55947 16652 55989 16661
rect 55947 16612 55948 16652
rect 55988 16612 55989 16652
rect 55947 16603 55989 16612
rect 55660 16232 55700 16603
rect 55756 16484 55796 16493
rect 56044 16484 56084 17032
rect 55796 16444 56084 16484
rect 55756 16435 55796 16444
rect 55660 16183 55700 16192
rect 56140 16232 56180 17116
rect 56455 17072 56495 17472
rect 56745 17240 56785 17472
rect 56236 17032 56495 17072
rect 56620 17200 56785 17240
rect 56236 16484 56276 17032
rect 56620 16988 56660 17200
rect 56855 17072 56895 17472
rect 57145 17156 57185 17472
rect 56236 16435 56276 16444
rect 56524 16948 56660 16988
rect 56812 17032 56895 17072
rect 57100 17116 57185 17156
rect 56524 16241 56564 16948
rect 56812 16736 56852 17032
rect 56620 16696 56852 16736
rect 56620 16484 56660 16696
rect 56620 16435 56660 16444
rect 55412 16108 55604 16148
rect 55372 16099 55412 16108
rect 56140 16073 56180 16192
rect 56523 16232 56565 16241
rect 56908 16232 56948 16241
rect 57100 16232 57140 17116
rect 57255 17072 57295 17472
rect 57545 17156 57585 17472
rect 56523 16192 56524 16232
rect 56564 16192 56565 16232
rect 56523 16183 56565 16192
rect 56812 16192 56908 16232
rect 56948 16192 57140 16232
rect 57196 17032 57295 17072
rect 57484 17116 57585 17156
rect 56139 16064 56181 16073
rect 56139 16024 56140 16064
rect 56180 16024 56181 16064
rect 56139 16015 56181 16024
rect 55467 15980 55509 15989
rect 55467 15940 55468 15980
rect 55508 15940 55509 15980
rect 55467 15931 55509 15940
rect 54603 15812 54645 15821
rect 54603 15772 54604 15812
rect 54644 15772 54645 15812
rect 54603 15763 54645 15772
rect 53643 15644 53685 15653
rect 53643 15604 53644 15644
rect 53684 15604 53685 15644
rect 53643 15595 53685 15604
rect 53548 15511 53588 15520
rect 53644 14048 53684 15595
rect 54412 15560 54452 15569
rect 54316 14888 54356 14897
rect 53067 13880 53109 13889
rect 53067 13840 53068 13880
rect 53108 13840 53109 13880
rect 53067 13831 53109 13840
rect 53452 13469 53492 14008
rect 53548 14008 53644 14048
rect 53548 13637 53588 14008
rect 53644 13999 53684 14008
rect 53835 14048 53877 14057
rect 53835 14008 53836 14048
rect 53876 14008 53877 14048
rect 53835 13999 53877 14008
rect 54220 14048 54260 14057
rect 54316 14048 54356 14848
rect 54412 14477 54452 15520
rect 54411 14468 54453 14477
rect 54411 14428 54412 14468
rect 54452 14428 54453 14468
rect 54411 14419 54453 14428
rect 54260 14008 54356 14048
rect 54220 13999 54260 14008
rect 53836 13914 53876 13999
rect 53644 13796 53684 13805
rect 53684 13756 54452 13796
rect 53644 13747 53684 13756
rect 53547 13628 53589 13637
rect 53547 13588 53548 13628
rect 53588 13588 53589 13628
rect 53547 13579 53589 13588
rect 53451 13460 53493 13469
rect 53451 13420 53452 13460
rect 53492 13420 53493 13460
rect 53451 13411 53493 13420
rect 53259 13208 53301 13217
rect 53259 13168 53260 13208
rect 53300 13168 53301 13208
rect 53259 13159 53301 13168
rect 54412 13208 54452 13756
rect 54507 13712 54549 13721
rect 54507 13672 54508 13712
rect 54548 13672 54549 13712
rect 54507 13663 54549 13672
rect 54412 13159 54452 13168
rect 54508 13208 54548 13663
rect 54508 13159 54548 13168
rect 51916 12940 52148 12980
rect 52588 12940 52820 12980
rect 51915 12872 51957 12881
rect 51915 12832 51916 12872
rect 51956 12832 51957 12872
rect 51915 12823 51957 12832
rect 51819 12704 51861 12713
rect 51819 12664 51820 12704
rect 51860 12664 51861 12704
rect 51819 12655 51861 12664
rect 51628 12487 51668 12496
rect 51819 12536 51861 12545
rect 51819 12496 51820 12536
rect 51860 12496 51861 12536
rect 51819 12487 51861 12496
rect 50763 11948 50805 11957
rect 50763 11908 50764 11948
rect 50804 11908 50805 11948
rect 50763 11899 50805 11908
rect 50379 11780 50421 11789
rect 50188 11740 50324 11780
rect 50284 11696 50324 11740
rect 50379 11740 50380 11780
rect 50420 11740 50421 11780
rect 50379 11731 50421 11740
rect 50188 11675 50228 11684
rect 50188 11621 50228 11635
rect 50187 11612 50229 11621
rect 50187 11572 50188 11612
rect 50228 11572 50229 11612
rect 50187 11563 50229 11572
rect 50188 11540 50228 11563
rect 49995 11024 50037 11033
rect 49995 10984 49996 11024
rect 50036 10984 50037 11024
rect 49995 10975 50037 10984
rect 50284 10361 50324 11656
rect 50380 11696 50420 11731
rect 50380 11646 50420 11656
rect 50764 11696 50804 11899
rect 50956 11696 50996 12487
rect 51820 12402 51860 12487
rect 51724 12284 51764 12293
rect 51628 12244 51724 12284
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 51436 11864 51476 11873
rect 51052 11696 51092 11705
rect 50956 11656 51052 11696
rect 50764 11647 50804 11656
rect 51052 11647 51092 11656
rect 51147 11612 51189 11621
rect 51147 11572 51148 11612
rect 51188 11572 51189 11612
rect 51147 11563 51189 11572
rect 50379 11528 50421 11537
rect 50379 11488 50380 11528
rect 50420 11488 50421 11528
rect 50379 11479 50421 11488
rect 50476 11528 50516 11537
rect 50516 11488 50804 11528
rect 50476 11479 50516 11488
rect 50380 11192 50420 11479
rect 50476 11192 50516 11201
rect 50380 11152 50476 11192
rect 50476 11143 50516 11152
rect 50764 11024 50804 11488
rect 51148 11478 51188 11563
rect 50956 11152 51284 11192
rect 50859 11108 50901 11117
rect 50859 11068 50860 11108
rect 50900 11068 50901 11108
rect 50859 11059 50901 11068
rect 50764 10975 50804 10984
rect 50860 10974 50900 11059
rect 50956 11024 50996 11152
rect 50956 10975 50996 10984
rect 51052 11024 51092 11033
rect 51052 10772 51092 10984
rect 51244 10856 51284 11152
rect 51340 11033 51380 11118
rect 51339 11024 51381 11033
rect 51339 10984 51340 11024
rect 51380 10984 51381 11024
rect 51436 11024 51476 11824
rect 51628 11696 51668 12244
rect 51724 12235 51764 12244
rect 51819 12116 51861 12125
rect 51819 12076 51820 12116
rect 51860 12076 51861 12116
rect 51819 12067 51861 12076
rect 51628 11647 51668 11656
rect 51724 11696 51764 11705
rect 51532 11024 51572 11033
rect 51436 10984 51532 11024
rect 51339 10975 51381 10984
rect 51532 10975 51572 10984
rect 51724 10940 51764 11656
rect 51820 11612 51860 12067
rect 51916 11948 51956 12823
rect 52012 12536 52052 12545
rect 52012 12125 52052 12496
rect 52011 12116 52053 12125
rect 52011 12076 52012 12116
rect 52052 12076 52053 12116
rect 52011 12067 52053 12076
rect 51916 11908 52052 11948
rect 51915 11696 51957 11705
rect 51915 11656 51916 11696
rect 51956 11656 51957 11696
rect 51915 11647 51957 11656
rect 51820 11563 51860 11572
rect 51916 11562 51956 11647
rect 51628 10900 51764 10940
rect 51916 10940 51956 10949
rect 52012 10940 52052 11908
rect 52108 11705 52148 12940
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 52396 12536 52436 12545
rect 52436 12496 52532 12536
rect 52396 12487 52436 12496
rect 52203 11864 52245 11873
rect 52203 11824 52204 11864
rect 52244 11824 52245 11864
rect 52203 11815 52245 11824
rect 52492 11864 52532 12496
rect 52492 11815 52532 11824
rect 52107 11696 52149 11705
rect 52107 11656 52108 11696
rect 52148 11656 52149 11696
rect 52107 11647 52149 11656
rect 52107 11528 52149 11537
rect 52107 11488 52108 11528
rect 52148 11488 52149 11528
rect 52107 11479 52149 11488
rect 51956 10900 52052 10940
rect 51436 10856 51476 10865
rect 51628 10856 51668 10900
rect 51916 10891 51956 10900
rect 51244 10816 51436 10856
rect 51476 10816 51668 10856
rect 51436 10807 51476 10816
rect 50956 10732 51092 10772
rect 51724 10772 51764 10781
rect 51764 10732 51860 10772
rect 50667 10688 50709 10697
rect 50667 10648 50668 10688
rect 50708 10648 50709 10688
rect 50667 10639 50709 10648
rect 50283 10352 50325 10361
rect 50283 10312 50284 10352
rect 50324 10312 50325 10352
rect 50283 10303 50325 10312
rect 50284 10184 50324 10193
rect 50324 10144 50420 10184
rect 50284 10135 50324 10144
rect 49900 10100 49940 10109
rect 49900 9689 49940 10060
rect 49899 9680 49941 9689
rect 49899 9640 49900 9680
rect 49940 9640 49941 9680
rect 49899 9631 49941 9640
rect 50380 9344 50420 10144
rect 50668 9512 50708 10639
rect 50668 9463 50708 9472
rect 49804 9304 50036 9344
rect 49899 9176 49941 9185
rect 49899 9136 49900 9176
rect 49940 9136 49941 9176
rect 49899 9127 49941 9136
rect 49227 8840 49269 8849
rect 49227 8800 49228 8840
rect 49268 8800 49269 8840
rect 49227 8791 49269 8800
rect 49324 8840 49364 8849
rect 48844 8345 48884 8632
rect 49036 8672 49076 8683
rect 49036 8597 49076 8632
rect 49131 8672 49173 8681
rect 49131 8632 49132 8672
rect 49172 8632 49173 8672
rect 49131 8623 49173 8632
rect 49035 8588 49077 8597
rect 49035 8548 49036 8588
rect 49076 8548 49077 8588
rect 49035 8539 49077 8548
rect 49132 8538 49172 8623
rect 48940 8504 48980 8513
rect 48843 8336 48885 8345
rect 48843 8296 48844 8336
rect 48884 8296 48885 8336
rect 48843 8287 48885 8296
rect 48940 8177 48980 8464
rect 48939 8168 48981 8177
rect 48939 8128 48940 8168
rect 48980 8128 48981 8168
rect 48939 8119 48981 8128
rect 48844 8009 48884 8094
rect 49228 8009 49268 8791
rect 48843 8000 48885 8009
rect 48843 7959 48844 8000
rect 48884 7959 48885 8000
rect 48843 7951 48885 7959
rect 49227 8000 49269 8009
rect 49227 7960 49228 8000
rect 49268 7960 49269 8000
rect 49227 7951 49269 7960
rect 48844 7950 48884 7951
rect 49228 7866 49268 7951
rect 48652 7783 48692 7792
rect 48747 7832 48789 7841
rect 48747 7792 48748 7832
rect 48788 7792 48789 7832
rect 48747 7783 48789 7792
rect 48460 7624 48692 7664
rect 48363 7412 48405 7421
rect 48363 7372 48364 7412
rect 48404 7372 48405 7412
rect 48363 7363 48405 7372
rect 48364 6488 48404 6497
rect 48172 6448 48364 6488
rect 48364 6439 48404 6448
rect 48556 6488 48596 6497
rect 48460 6236 48500 6245
rect 48460 5741 48500 6196
rect 48556 5909 48596 6448
rect 48555 5900 48597 5909
rect 48555 5860 48556 5900
rect 48596 5860 48597 5900
rect 48555 5851 48597 5860
rect 48459 5732 48501 5741
rect 48459 5692 48460 5732
rect 48500 5692 48501 5732
rect 48459 5683 48501 5692
rect 48076 5599 48116 5608
rect 48364 5648 48404 5659
rect 48364 5573 48404 5608
rect 48363 5564 48405 5573
rect 48268 5524 48364 5564
rect 48404 5524 48405 5564
rect 47883 5480 47925 5489
rect 47883 5440 47884 5480
rect 47924 5440 47925 5480
rect 47883 5431 47925 5440
rect 48268 4985 48308 5524
rect 48363 5515 48405 5524
rect 48460 5564 48500 5573
rect 48460 5144 48500 5524
rect 48364 5104 48500 5144
rect 48267 4976 48309 4985
rect 48267 4936 48268 4976
rect 48308 4936 48309 4976
rect 48267 4927 48309 4936
rect 48076 4724 48116 4733
rect 48076 4556 48116 4684
rect 48364 4556 48404 5104
rect 48555 5060 48597 5069
rect 48555 5020 48556 5060
rect 48596 5020 48597 5060
rect 48555 5011 48597 5020
rect 48459 4976 48501 4985
rect 48459 4936 48460 4976
rect 48500 4936 48501 4976
rect 48459 4927 48501 4936
rect 48460 4842 48500 4927
rect 48556 4926 48596 5011
rect 48652 4976 48692 7624
rect 48748 7160 48788 7783
rect 49035 7664 49077 7673
rect 49035 7624 49036 7664
rect 49076 7624 49077 7664
rect 49035 7615 49077 7624
rect 48748 7111 48788 7120
rect 48844 6488 48884 6497
rect 48747 5900 48789 5909
rect 48747 5860 48748 5900
rect 48788 5860 48789 5900
rect 48844 5900 48884 6448
rect 48940 5900 48980 5909
rect 48844 5860 48940 5900
rect 48747 5851 48789 5860
rect 48940 5851 48980 5860
rect 48748 5766 48788 5851
rect 48940 5648 48980 5657
rect 49036 5648 49076 7615
rect 49132 7160 49172 7169
rect 49324 7160 49364 8800
rect 49708 8672 49748 8681
rect 49708 7757 49748 8632
rect 49803 8672 49845 8681
rect 49803 8632 49804 8672
rect 49844 8632 49845 8672
rect 49803 8623 49845 8632
rect 49900 8672 49940 9127
rect 49996 8681 50036 9304
rect 50380 9295 50420 9304
rect 50763 9176 50805 9185
rect 50763 9136 50764 9176
rect 50804 9136 50805 9176
rect 50763 9127 50805 9136
rect 49804 8538 49844 8623
rect 49900 8261 49940 8632
rect 49995 8672 50037 8681
rect 49995 8632 49996 8672
rect 50036 8632 50037 8672
rect 49995 8623 50037 8632
rect 50187 8588 50229 8597
rect 50187 8548 50188 8588
rect 50228 8548 50229 8588
rect 50187 8539 50229 8548
rect 49899 8252 49941 8261
rect 49899 8212 49900 8252
rect 49940 8212 49941 8252
rect 49899 8203 49941 8212
rect 50188 8000 50228 8539
rect 50188 7951 50228 7960
rect 50476 8000 50516 8009
rect 49707 7748 49749 7757
rect 49707 7708 49708 7748
rect 49748 7708 49749 7748
rect 49707 7699 49749 7708
rect 49900 7748 49940 7757
rect 49940 7708 50036 7748
rect 49900 7699 49940 7708
rect 49172 7120 49364 7160
rect 49996 7160 50036 7708
rect 50476 7253 50516 7960
rect 50764 7496 50804 9127
rect 50956 8924 50996 10732
rect 51724 10723 51764 10732
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 51148 10184 51188 10193
rect 51188 10144 51764 10184
rect 51148 10135 51188 10144
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 51340 8924 51380 8933
rect 50956 8884 51340 8924
rect 51340 8875 51380 8884
rect 51531 8840 51573 8849
rect 50956 8798 50996 8807
rect 51531 8800 51532 8840
rect 51572 8800 51573 8840
rect 51531 8791 51573 8800
rect 50860 8000 50900 8009
rect 50956 8000 50996 8758
rect 51339 8672 51381 8681
rect 51339 8632 51340 8672
rect 51380 8632 51381 8672
rect 51339 8623 51381 8632
rect 51532 8672 51572 8791
rect 51627 8756 51669 8765
rect 51627 8716 51628 8756
rect 51668 8716 51669 8756
rect 51627 8707 51669 8716
rect 51532 8623 51572 8632
rect 51628 8672 51668 8707
rect 51340 8538 51380 8623
rect 51628 8621 51668 8632
rect 51724 8513 51764 10144
rect 51820 8849 51860 10732
rect 52011 10352 52053 10361
rect 52011 10312 52012 10352
rect 52052 10312 52053 10352
rect 52011 10303 52053 10312
rect 51915 8924 51957 8933
rect 51915 8884 51916 8924
rect 51956 8884 51957 8924
rect 51915 8875 51957 8884
rect 51819 8840 51861 8849
rect 51819 8800 51820 8840
rect 51860 8800 51861 8840
rect 51819 8791 51861 8800
rect 51723 8504 51765 8513
rect 51723 8464 51724 8504
rect 51764 8464 51765 8504
rect 51723 8455 51765 8464
rect 50900 7960 50996 8000
rect 51724 8000 51764 8455
rect 50860 7951 50900 7960
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 50764 7456 50996 7496
rect 50956 7412 50996 7456
rect 51148 7412 51188 7421
rect 50956 7372 51148 7412
rect 51148 7363 51188 7372
rect 50475 7244 50517 7253
rect 50475 7204 50476 7244
rect 50516 7204 50517 7244
rect 50475 7195 50517 7204
rect 50036 7120 50132 7160
rect 49132 7111 49172 7120
rect 49996 7111 50036 7120
rect 50092 6497 50132 7120
rect 51724 6497 51764 7960
rect 51916 7496 51956 8875
rect 52012 8504 52052 10303
rect 52108 9605 52148 11479
rect 52204 11192 52244 11815
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 52204 11152 52724 11192
rect 52684 10184 52724 11152
rect 52300 10025 52340 10110
rect 52684 10025 52724 10144
rect 52299 10016 52341 10025
rect 52204 9976 52300 10016
rect 52340 9976 52341 10016
rect 52107 9596 52149 9605
rect 52107 9556 52108 9596
rect 52148 9556 52149 9596
rect 52107 9547 52149 9556
rect 52108 9428 52148 9437
rect 52108 8681 52148 9388
rect 52204 8765 52244 9976
rect 52299 9967 52341 9976
rect 52683 10016 52725 10025
rect 52683 9976 52684 10016
rect 52724 9976 52725 10016
rect 52683 9967 52725 9976
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 52684 9680 52724 9689
rect 52780 9680 52820 12940
rect 53260 12536 53300 13159
rect 54604 13049 54644 15763
rect 55083 14468 55125 14477
rect 55083 14428 55084 14468
rect 55124 14428 55125 14468
rect 55083 14419 55125 14428
rect 54699 14048 54741 14057
rect 54699 14008 54700 14048
rect 54740 14008 54741 14048
rect 54699 13999 54741 14008
rect 55084 14048 55124 14419
rect 55084 13999 55124 14008
rect 54700 13460 54740 13999
rect 54700 13411 54740 13420
rect 55179 13292 55221 13301
rect 55179 13252 55180 13292
rect 55220 13252 55221 13292
rect 55179 13243 55221 13252
rect 54700 13208 54740 13217
rect 55084 13208 55124 13217
rect 54740 13168 55084 13208
rect 54700 13159 54740 13168
rect 55084 13159 55124 13168
rect 55180 13208 55220 13243
rect 55180 13157 55220 13168
rect 55276 13208 55316 13219
rect 55276 13133 55316 13168
rect 55371 13208 55413 13217
rect 55371 13168 55372 13208
rect 55412 13168 55413 13208
rect 55371 13159 55413 13168
rect 55275 13124 55317 13133
rect 55275 13084 55276 13124
rect 55316 13084 55317 13124
rect 55275 13075 55317 13084
rect 55372 13074 55412 13159
rect 54603 13040 54645 13049
rect 54603 13000 54604 13040
rect 54644 13000 54645 13040
rect 54603 12991 54645 13000
rect 54891 13040 54933 13049
rect 54891 13000 54892 13040
rect 54932 13000 54933 13040
rect 54891 12991 54933 13000
rect 54892 12620 54932 12991
rect 54892 12571 54932 12580
rect 55468 12545 55508 15931
rect 55563 15476 55605 15485
rect 55563 15436 55564 15476
rect 55604 15436 55605 15476
rect 55563 15427 55605 15436
rect 55564 15317 55604 15427
rect 55563 15308 55605 15317
rect 55563 15268 55564 15308
rect 55604 15268 55605 15308
rect 55563 15259 55605 15268
rect 56716 14888 56756 14897
rect 56620 14848 56716 14888
rect 56043 14720 56085 14729
rect 56043 14680 56044 14720
rect 56084 14680 56085 14720
rect 56043 14671 56085 14680
rect 56331 14720 56373 14729
rect 56331 14680 56332 14720
rect 56372 14680 56373 14720
rect 56331 14671 56373 14680
rect 56044 14586 56084 14671
rect 56332 14586 56372 14671
rect 56428 14636 56468 14645
rect 55947 14468 55989 14477
rect 55947 14428 55948 14468
rect 55988 14428 55989 14468
rect 55947 14419 55989 14428
rect 55948 12980 55988 14419
rect 56428 14300 56468 14596
rect 56236 14260 56468 14300
rect 56236 14216 56276 14260
rect 56236 14167 56276 14176
rect 56428 14048 56468 14057
rect 56428 13889 56468 14008
rect 56620 14048 56660 14848
rect 56716 14839 56756 14848
rect 56620 13999 56660 14008
rect 56427 13880 56469 13889
rect 56427 13840 56428 13880
rect 56468 13840 56469 13880
rect 56427 13831 56469 13840
rect 56236 13796 56276 13805
rect 56044 13756 56236 13796
rect 56044 13217 56084 13756
rect 56236 13747 56276 13756
rect 56524 13796 56564 13807
rect 56524 13721 56564 13756
rect 56523 13712 56565 13721
rect 56523 13672 56524 13712
rect 56564 13672 56565 13712
rect 56523 13663 56565 13672
rect 56235 13628 56277 13637
rect 56235 13588 56236 13628
rect 56276 13588 56277 13628
rect 56235 13579 56277 13588
rect 56139 13460 56181 13469
rect 56139 13420 56140 13460
rect 56180 13420 56181 13460
rect 56139 13411 56181 13420
rect 56043 13208 56085 13217
rect 56043 13168 56044 13208
rect 56084 13168 56085 13208
rect 56043 13159 56085 13168
rect 56140 13208 56180 13411
rect 56236 13208 56276 13579
rect 56812 13553 56852 16192
rect 56908 16183 56948 16192
rect 57004 16064 57044 16073
rect 57196 16064 57236 17032
rect 57484 16988 57524 17116
rect 57655 17072 57695 17472
rect 57945 17165 57985 17472
rect 57944 17156 57986 17165
rect 57944 17116 57945 17156
rect 57985 17116 58004 17156
rect 57944 17107 58004 17116
rect 57292 16948 57524 16988
rect 57580 17032 57695 17072
rect 57292 16493 57332 16948
rect 57580 16568 57620 17032
rect 57388 16528 57620 16568
rect 57291 16484 57333 16493
rect 57291 16444 57292 16484
rect 57332 16444 57333 16484
rect 57291 16435 57333 16444
rect 57388 16484 57428 16528
rect 57388 16435 57428 16444
rect 57292 16232 57332 16435
rect 57580 16400 57620 16409
rect 57292 16183 57332 16192
rect 57484 16360 57580 16400
rect 57044 16024 57236 16064
rect 57291 16064 57333 16073
rect 57291 16024 57292 16064
rect 57332 16024 57333 16064
rect 57004 16015 57044 16024
rect 57291 16015 57333 16024
rect 57100 15560 57140 15569
rect 56908 15520 57100 15560
rect 56908 14972 56948 15520
rect 57100 15511 57140 15520
rect 57003 15308 57045 15317
rect 57003 15268 57004 15308
rect 57044 15268 57045 15308
rect 57003 15259 57045 15268
rect 56908 14923 56948 14932
rect 56908 14720 56948 14729
rect 56908 14561 56948 14680
rect 56907 14552 56949 14561
rect 56907 14512 56908 14552
rect 56948 14512 56949 14552
rect 56907 14503 56949 14512
rect 56811 13544 56853 13553
rect 56811 13504 56812 13544
rect 56852 13504 56853 13544
rect 56811 13495 56853 13504
rect 56332 13376 56372 13385
rect 56372 13336 56852 13376
rect 56332 13327 56372 13336
rect 56331 13208 56373 13217
rect 56236 13168 56332 13208
rect 56372 13168 56373 13208
rect 56140 13159 56180 13168
rect 56331 13159 56373 13168
rect 56524 13208 56564 13217
rect 56332 13074 56372 13159
rect 56427 13124 56469 13133
rect 56427 13084 56428 13124
rect 56468 13084 56469 13124
rect 56427 13075 56469 13084
rect 55948 12940 56180 12980
rect 56140 12545 56180 12940
rect 53260 12487 53300 12496
rect 54411 12536 54453 12545
rect 54411 12496 54412 12536
rect 54452 12496 54453 12536
rect 54411 12487 54453 12496
rect 55276 12536 55316 12545
rect 54412 12452 54452 12487
rect 54412 12401 54452 12412
rect 55276 11864 55316 12496
rect 55467 12536 55509 12545
rect 55467 12496 55468 12536
rect 55508 12496 55509 12536
rect 55467 12487 55509 12496
rect 56139 12536 56181 12545
rect 56139 12496 56140 12536
rect 56180 12496 56181 12536
rect 56139 12487 56181 12496
rect 56140 12402 56180 12487
rect 56235 12200 56277 12209
rect 56235 12160 56236 12200
rect 56276 12160 56277 12200
rect 56235 12151 56277 12160
rect 55372 11864 55412 11873
rect 53740 11824 54068 11864
rect 55276 11824 55372 11864
rect 53355 11696 53397 11705
rect 53355 11656 53356 11696
rect 53396 11656 53397 11696
rect 53355 11647 53397 11656
rect 53740 11696 53780 11824
rect 53740 11647 53780 11656
rect 53931 11696 53973 11705
rect 53931 11656 53932 11696
rect 53972 11656 53973 11696
rect 53931 11647 53973 11656
rect 53356 11033 53396 11647
rect 53836 11612 53876 11621
rect 53836 11276 53876 11572
rect 53644 11236 53876 11276
rect 53355 11024 53397 11033
rect 53355 10984 53356 11024
rect 53396 10984 53397 11024
rect 53355 10975 53397 10984
rect 53548 11024 53588 11033
rect 53356 10890 53396 10975
rect 53355 10772 53397 10781
rect 53355 10732 53356 10772
rect 53396 10732 53397 10772
rect 53548 10772 53588 10984
rect 53644 11024 53684 11236
rect 53739 11108 53781 11117
rect 53739 11068 53740 11108
rect 53780 11068 53781 11108
rect 53739 11059 53781 11068
rect 53644 10975 53684 10984
rect 53548 10732 53684 10772
rect 53355 10723 53397 10732
rect 53356 10638 53396 10723
rect 53356 10352 53396 10361
rect 53396 10312 53588 10352
rect 53356 10303 53396 10312
rect 52971 10184 53013 10193
rect 52971 10144 52972 10184
rect 53012 10144 53013 10184
rect 52971 10135 53013 10144
rect 53548 10184 53588 10312
rect 53548 10135 53588 10144
rect 52972 10050 53012 10135
rect 53644 10109 53684 10732
rect 53740 10184 53780 11059
rect 53836 11024 53876 11033
rect 53836 10781 53876 10984
rect 53835 10772 53877 10781
rect 53835 10732 53836 10772
rect 53876 10732 53877 10772
rect 53835 10723 53877 10732
rect 53932 10193 53972 11647
rect 53068 10100 53108 10109
rect 53068 9941 53108 10060
rect 53163 10100 53205 10109
rect 53163 10060 53164 10100
rect 53204 10060 53205 10100
rect 53163 10051 53205 10060
rect 53643 10100 53685 10109
rect 53643 10060 53644 10100
rect 53684 10060 53685 10100
rect 53643 10051 53685 10060
rect 53067 9932 53109 9941
rect 53067 9892 53068 9932
rect 53108 9892 53109 9932
rect 53067 9883 53109 9892
rect 52724 9640 52820 9680
rect 53067 9680 53109 9689
rect 53067 9640 53068 9680
rect 53108 9640 53109 9680
rect 52684 9631 52724 9640
rect 53067 9631 53109 9640
rect 52395 9596 52437 9605
rect 52395 9556 52396 9596
rect 52436 9556 52437 9596
rect 52395 9547 52437 9556
rect 52203 8756 52245 8765
rect 52203 8716 52204 8756
rect 52244 8716 52245 8756
rect 52203 8707 52245 8716
rect 52107 8672 52149 8681
rect 52107 8632 52108 8672
rect 52148 8632 52149 8672
rect 52107 8623 52149 8632
rect 52204 8672 52244 8707
rect 52396 8681 52436 9547
rect 53068 9546 53108 9631
rect 52972 9512 53012 9521
rect 52492 9472 52972 9512
rect 52204 8622 52244 8632
rect 52300 8672 52340 8681
rect 52300 8504 52340 8632
rect 52395 8672 52437 8681
rect 52395 8632 52396 8672
rect 52436 8632 52437 8672
rect 52395 8623 52437 8632
rect 52492 8672 52532 9472
rect 52972 9463 53012 9472
rect 53164 9512 53204 10051
rect 53451 10016 53493 10025
rect 53451 9976 53452 10016
rect 53492 9976 53493 10016
rect 53451 9967 53493 9976
rect 53164 9463 53204 9472
rect 53270 9493 53310 9502
rect 52683 9260 52725 9269
rect 52683 9220 52684 9260
rect 52724 9220 52725 9260
rect 52683 9211 52725 9220
rect 52684 9126 52724 9211
rect 53270 9092 53310 9453
rect 53270 9052 53396 9092
rect 52683 8924 52725 8933
rect 52683 8884 52684 8924
rect 52724 8884 52725 8924
rect 52683 8875 52725 8884
rect 53259 8924 53301 8933
rect 53259 8884 53260 8924
rect 53300 8884 53301 8924
rect 53259 8875 53301 8884
rect 52492 8623 52532 8632
rect 52684 8672 52724 8875
rect 52875 8840 52917 8849
rect 52875 8800 52876 8840
rect 52916 8800 52917 8840
rect 52875 8791 52917 8800
rect 52684 8623 52724 8632
rect 52876 8672 52916 8791
rect 53260 8689 53300 8875
rect 52876 8623 52916 8632
rect 52972 8672 53012 8681
rect 52396 8538 52436 8623
rect 52012 8464 52340 8504
rect 52779 8504 52821 8513
rect 52779 8464 52780 8504
rect 52820 8464 52821 8504
rect 52204 8093 52244 8464
rect 52779 8455 52821 8464
rect 52780 8370 52820 8455
rect 52972 8429 53012 8632
rect 53163 8672 53205 8681
rect 53163 8632 53164 8672
rect 53204 8632 53205 8672
rect 53260 8640 53300 8649
rect 53163 8623 53205 8632
rect 52971 8420 53013 8429
rect 52971 8380 52972 8420
rect 53012 8380 53013 8420
rect 52971 8371 53013 8380
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 52876 8168 52916 8177
rect 52972 8168 53012 8371
rect 52916 8128 53012 8168
rect 52876 8119 52916 8128
rect 52203 8084 52245 8093
rect 52203 8044 52204 8084
rect 52244 8044 52245 8084
rect 52203 8035 52245 8044
rect 52683 8084 52725 8093
rect 52683 8044 52684 8084
rect 52724 8044 52725 8084
rect 52683 8035 52725 8044
rect 51916 7456 52052 7496
rect 51916 7328 51956 7337
rect 49228 6488 49268 6497
rect 49228 5816 49268 6448
rect 50091 6488 50133 6497
rect 50091 6448 50092 6488
rect 50132 6448 50133 6488
rect 50091 6439 50133 6448
rect 50859 6488 50901 6497
rect 50859 6448 50860 6488
rect 50900 6448 50901 6488
rect 50859 6439 50901 6448
rect 51436 6488 51476 6497
rect 50092 6354 50132 6439
rect 50379 6152 50421 6161
rect 50379 6112 50380 6152
rect 50420 6112 50421 6152
rect 50379 6103 50421 6112
rect 49420 5816 49460 5825
rect 49228 5776 49420 5816
rect 49420 5767 49460 5776
rect 48980 5608 49076 5648
rect 49131 5648 49173 5657
rect 49131 5608 49132 5648
rect 49172 5608 49173 5648
rect 48940 5599 48980 5608
rect 49131 5599 49173 5608
rect 49228 5648 49268 5657
rect 49132 5514 49172 5599
rect 48939 5480 48981 5489
rect 48939 5440 48940 5480
rect 48980 5440 48981 5480
rect 48939 5431 48981 5440
rect 48652 4927 48692 4936
rect 48844 4976 48884 4985
rect 48844 4556 48884 4936
rect 48940 4976 48980 5431
rect 49131 5144 49173 5153
rect 49131 5104 49132 5144
rect 49172 5104 49173 5144
rect 49131 5095 49173 5104
rect 48940 4927 48980 4936
rect 49132 4976 49172 5095
rect 49228 5069 49268 5608
rect 50380 5573 50420 6103
rect 50379 5564 50421 5573
rect 50379 5524 50380 5564
rect 50420 5524 50421 5564
rect 50379 5515 50421 5524
rect 49227 5060 49269 5069
rect 49227 5020 49228 5060
rect 49268 5020 49269 5060
rect 49227 5011 49269 5020
rect 49132 4927 49172 4936
rect 50092 4808 50132 4817
rect 49132 4724 49172 4733
rect 49172 4684 49940 4724
rect 49132 4675 49172 4684
rect 48076 4516 48884 4556
rect 47596 4087 47636 4096
rect 47692 4136 47732 4145
rect 48076 4136 48116 4516
rect 47732 4096 48116 4136
rect 47692 4087 47732 4096
rect 47116 3928 47540 3968
rect 49612 4052 49652 4061
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 49612 3641 49652 4012
rect 49611 3632 49653 3641
rect 49611 3592 49612 3632
rect 49652 3592 49653 3632
rect 49611 3583 49653 3592
rect 49900 3464 49940 4684
rect 49996 4136 50036 4145
rect 50092 4136 50132 4768
rect 50667 4220 50709 4229
rect 50667 4180 50668 4220
rect 50708 4180 50709 4220
rect 50667 4171 50709 4180
rect 50036 4096 50132 4136
rect 49996 4087 50036 4096
rect 50187 3632 50229 3641
rect 50187 3592 50188 3632
rect 50228 3592 50229 3632
rect 50187 3583 50229 3592
rect 50188 3498 50228 3583
rect 49996 3464 50036 3473
rect 49900 3424 49996 3464
rect 49996 3415 50036 3424
rect 50092 3464 50132 3473
rect 50092 3305 50132 3424
rect 50284 3464 50324 3473
rect 50572 3464 50612 3473
rect 50324 3424 50572 3464
rect 50284 3415 50324 3424
rect 50572 3415 50612 3424
rect 50668 3464 50708 4171
rect 50860 4136 50900 6439
rect 51244 6245 51284 6330
rect 51436 6245 51476 6448
rect 51723 6488 51765 6497
rect 51723 6448 51724 6488
rect 51764 6448 51765 6488
rect 51723 6439 51765 6448
rect 51820 6488 51860 6497
rect 51916 6488 51956 7288
rect 51860 6448 51956 6488
rect 51820 6439 51860 6448
rect 51243 6236 51285 6245
rect 51243 6196 51244 6236
rect 51284 6196 51285 6236
rect 51243 6187 51285 6196
rect 51435 6236 51477 6245
rect 51435 6196 51436 6236
rect 51476 6196 51477 6236
rect 51435 6187 51477 6196
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 52012 5153 52052 7456
rect 52684 6992 52724 8035
rect 53068 8000 53108 8009
rect 52780 7960 53068 8000
rect 52780 7160 52820 7960
rect 53068 7951 53108 7960
rect 53164 8000 53204 8623
rect 53356 8513 53396 9052
rect 53452 9017 53492 9967
rect 53644 9966 53684 10051
rect 53740 9521 53780 10144
rect 53931 10184 53973 10193
rect 53931 10144 53932 10184
rect 53972 10144 53973 10184
rect 53931 10135 53973 10144
rect 53739 9512 53781 9521
rect 53739 9472 53740 9512
rect 53780 9472 53781 9512
rect 53739 9463 53781 9472
rect 53932 9512 53972 9521
rect 53740 9378 53780 9463
rect 53836 9260 53876 9269
rect 53451 9008 53493 9017
rect 53451 8968 53452 9008
rect 53492 8968 53493 9008
rect 53451 8959 53493 8968
rect 53452 8681 53492 8959
rect 53547 8924 53589 8933
rect 53547 8884 53548 8924
rect 53588 8884 53589 8924
rect 53547 8875 53589 8884
rect 53451 8672 53493 8681
rect 53451 8632 53452 8672
rect 53492 8632 53493 8672
rect 53451 8623 53493 8632
rect 53548 8672 53588 8875
rect 53739 8840 53781 8849
rect 53739 8800 53740 8840
rect 53780 8800 53781 8840
rect 53739 8791 53781 8800
rect 53548 8623 53588 8632
rect 53644 8588 53684 8597
rect 53355 8504 53397 8513
rect 53355 8464 53356 8504
rect 53396 8464 53397 8504
rect 53355 8455 53397 8464
rect 53644 8429 53684 8548
rect 53643 8420 53685 8429
rect 53643 8380 53644 8420
rect 53684 8380 53685 8420
rect 53643 8371 53685 8380
rect 53259 8084 53301 8093
rect 53259 8044 53260 8084
rect 53300 8044 53301 8084
rect 53259 8035 53301 8044
rect 52971 7832 53013 7841
rect 52971 7792 52972 7832
rect 53012 7792 53013 7832
rect 52971 7783 53013 7792
rect 52875 7244 52917 7253
rect 52875 7204 52876 7244
rect 52916 7204 52917 7244
rect 52875 7195 52917 7204
rect 52780 7111 52820 7120
rect 52876 7076 52916 7195
rect 52972 7160 53012 7783
rect 52972 7111 53012 7120
rect 53067 7160 53109 7169
rect 53067 7120 53068 7160
rect 53108 7120 53109 7160
rect 53067 7111 53109 7120
rect 52876 7027 52916 7036
rect 53068 7026 53108 7111
rect 52684 6952 52820 6992
rect 52780 6908 52820 6952
rect 52780 6868 52916 6908
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 52684 6488 52724 6497
rect 52395 6236 52437 6245
rect 52395 6196 52396 6236
rect 52436 6196 52437 6236
rect 52395 6187 52437 6196
rect 52204 5648 52244 5657
rect 52011 5144 52053 5153
rect 52011 5104 52012 5144
rect 52052 5104 52053 5144
rect 52011 5095 52053 5104
rect 52204 5144 52244 5608
rect 52299 5648 52341 5657
rect 52299 5608 52300 5648
rect 52340 5608 52341 5648
rect 52299 5599 52341 5608
rect 52300 5514 52340 5599
rect 52396 5564 52436 6187
rect 52684 5741 52724 6448
rect 52779 5816 52821 5825
rect 52779 5776 52780 5816
rect 52820 5776 52821 5816
rect 52779 5767 52821 5776
rect 52683 5732 52725 5741
rect 52683 5692 52684 5732
rect 52724 5692 52725 5732
rect 52683 5683 52725 5692
rect 52492 5648 52532 5657
rect 52780 5648 52820 5767
rect 52532 5608 52628 5648
rect 52492 5599 52532 5608
rect 52588 5564 52628 5608
rect 52780 5599 52820 5608
rect 52876 5648 52916 6868
rect 53164 5825 53204 7960
rect 53260 8021 53300 8035
rect 53260 7949 53300 7981
rect 53356 8000 53396 8009
rect 53644 8000 53684 8371
rect 53396 7960 53684 8000
rect 53356 7951 53396 7960
rect 53452 7253 53492 7284
rect 53740 7253 53780 8791
rect 53836 8009 53876 9220
rect 53932 8924 53972 9472
rect 53932 8875 53972 8884
rect 54028 8849 54068 11824
rect 55372 11815 55412 11824
rect 56236 11705 56276 12151
rect 56332 11864 56372 11873
rect 56235 11696 56277 11705
rect 56235 11656 56236 11696
rect 56276 11656 56277 11696
rect 56235 11647 56277 11656
rect 56236 11192 56276 11647
rect 56332 11444 56372 11824
rect 56428 11528 56468 13075
rect 56524 11696 56564 13168
rect 56715 13208 56757 13217
rect 56715 13168 56716 13208
rect 56756 13168 56757 13208
rect 56715 13159 56757 13168
rect 56812 13208 56852 13336
rect 56907 13292 56949 13301
rect 56907 13252 56908 13292
rect 56948 13252 56949 13292
rect 56907 13243 56949 13252
rect 56812 13159 56852 13168
rect 56620 13049 56660 13134
rect 56716 13074 56756 13159
rect 56619 13040 56661 13049
rect 56619 13000 56620 13040
rect 56660 13000 56661 13040
rect 56619 12991 56661 13000
rect 56908 12368 56948 13243
rect 56524 11647 56564 11656
rect 56620 12328 56948 12368
rect 56620 11696 56660 12328
rect 56811 11780 56853 11789
rect 56811 11740 56812 11780
rect 56852 11740 56853 11780
rect 56811 11731 56853 11740
rect 56620 11647 56660 11656
rect 56716 11696 56756 11705
rect 56716 11528 56756 11656
rect 56812 11696 56852 11731
rect 56812 11645 56852 11656
rect 56428 11488 56756 11528
rect 56332 11404 56852 11444
rect 56236 11143 56276 11152
rect 54123 11024 54165 11033
rect 54123 10984 54124 11024
rect 54164 10984 54165 11024
rect 54123 10975 54165 10984
rect 54220 11024 54260 11033
rect 55084 11024 55124 11033
rect 54260 10984 54356 11024
rect 54220 10975 54260 10984
rect 54027 8840 54069 8849
rect 54027 8800 54028 8840
rect 54068 8800 54069 8840
rect 54027 8791 54069 8800
rect 53931 8672 53973 8681
rect 54124 8672 54164 10975
rect 54316 10352 54356 10984
rect 54316 10303 54356 10312
rect 54220 9512 54260 9521
rect 54220 9017 54260 9472
rect 54412 9512 54452 9521
rect 54316 9260 54356 9269
rect 54219 9008 54261 9017
rect 54219 8968 54220 9008
rect 54260 8968 54261 9008
rect 54219 8959 54261 8968
rect 53931 8632 53932 8672
rect 53972 8632 53973 8672
rect 53931 8623 53973 8632
rect 54028 8632 54164 8672
rect 53835 8000 53877 8009
rect 53835 7960 53836 8000
rect 53876 7960 53877 8000
rect 53835 7951 53877 7960
rect 53451 7244 53493 7253
rect 53451 7204 53452 7244
rect 53492 7204 53493 7244
rect 53451 7195 53493 7204
rect 53739 7244 53781 7253
rect 53739 7204 53740 7244
rect 53780 7204 53781 7244
rect 53739 7195 53781 7204
rect 53452 7160 53492 7195
rect 53260 7118 53300 7127
rect 53260 6740 53300 7078
rect 53355 7076 53397 7085
rect 53355 7036 53356 7076
rect 53396 7036 53397 7076
rect 53355 7027 53397 7036
rect 53356 6942 53396 7027
rect 53260 6700 53396 6740
rect 53163 5816 53205 5825
rect 53068 5776 53164 5816
rect 53204 5776 53205 5816
rect 52684 5564 52724 5573
rect 52588 5524 52684 5564
rect 52396 5515 52436 5524
rect 52684 5515 52724 5524
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 52204 5095 52244 5104
rect 52299 5144 52341 5153
rect 52299 5104 52300 5144
rect 52340 5104 52341 5144
rect 52299 5095 52341 5104
rect 51819 5060 51861 5069
rect 51819 5020 51820 5060
rect 51860 5020 51861 5060
rect 51819 5011 51861 5020
rect 51532 4976 51572 4985
rect 51724 4976 51764 4985
rect 51572 4936 51668 4976
rect 51532 4927 51572 4936
rect 51628 4817 51668 4936
rect 51627 4808 51669 4817
rect 51627 4768 51628 4808
rect 51668 4768 51669 4808
rect 51627 4759 51669 4768
rect 51532 4724 51572 4733
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 51532 4397 51572 4684
rect 51531 4388 51573 4397
rect 51531 4348 51532 4388
rect 51572 4348 51573 4388
rect 51531 4339 51573 4348
rect 50860 4061 50900 4096
rect 50859 4052 50901 4061
rect 50859 4012 50860 4052
rect 50900 4012 50901 4052
rect 50859 4003 50901 4012
rect 50763 3968 50805 3977
rect 50763 3928 50764 3968
rect 50804 3928 50805 3968
rect 50763 3919 50805 3928
rect 50668 3415 50708 3424
rect 50764 3464 50804 3919
rect 50859 3632 50901 3641
rect 50859 3592 50860 3632
rect 50900 3592 50901 3632
rect 50859 3583 50901 3592
rect 50764 3415 50804 3424
rect 50860 3464 50900 3583
rect 50860 3415 50900 3424
rect 51627 3464 51669 3473
rect 51627 3424 51628 3464
rect 51668 3424 51669 3464
rect 51627 3415 51669 3424
rect 51628 3330 51668 3415
rect 51724 3305 51764 4936
rect 51820 4976 51860 5011
rect 51820 4925 51860 4936
rect 52012 4976 52052 4985
rect 52012 4388 52052 4936
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 52300 4976 52340 5095
rect 52587 5060 52629 5069
rect 52587 5020 52588 5060
rect 52628 5020 52629 5060
rect 52587 5011 52629 5020
rect 52300 4927 52340 4936
rect 52491 4976 52533 4985
rect 52491 4936 52492 4976
rect 52532 4936 52533 4976
rect 52491 4927 52533 4936
rect 52108 4842 52148 4927
rect 52492 4842 52532 4927
rect 52588 4926 52628 5011
rect 52684 4976 52724 4985
rect 52876 4976 52916 5608
rect 52971 5648 53013 5657
rect 52971 5608 52972 5648
rect 53012 5608 53013 5648
rect 52971 5599 53013 5608
rect 52972 5514 53012 5599
rect 52876 4936 53012 4976
rect 52012 4339 52052 4348
rect 52299 4388 52341 4397
rect 52299 4348 52300 4388
rect 52340 4348 52341 4388
rect 52299 4339 52341 4348
rect 51915 4304 51957 4313
rect 51915 4264 51916 4304
rect 51956 4264 51957 4304
rect 51915 4255 51957 4264
rect 51916 3464 51956 4255
rect 52300 4136 52340 4339
rect 52684 4313 52724 4936
rect 52876 4808 52916 4817
rect 52683 4304 52725 4313
rect 52683 4264 52684 4304
rect 52724 4264 52725 4304
rect 52683 4255 52725 4264
rect 52300 4087 52340 4096
rect 52684 4136 52724 4145
rect 52876 4136 52916 4768
rect 52724 4096 52916 4136
rect 52684 4087 52724 4096
rect 52972 3977 53012 4936
rect 53068 4229 53108 5776
rect 53163 5767 53205 5776
rect 53259 5060 53301 5069
rect 53356 5060 53396 6700
rect 53164 5020 53260 5060
rect 53300 5020 53396 5060
rect 53067 4220 53109 4229
rect 53067 4180 53068 4220
rect 53108 4180 53109 4220
rect 53067 4171 53109 4180
rect 52012 3968 52052 3977
rect 52012 3641 52052 3928
rect 52971 3968 53013 3977
rect 52971 3928 52972 3968
rect 53012 3928 53013 3968
rect 52971 3919 53013 3928
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 52011 3632 52053 3641
rect 52011 3592 52012 3632
rect 52052 3592 52053 3632
rect 52011 3583 52053 3592
rect 52012 3548 52052 3583
rect 52012 3497 52052 3508
rect 51916 3415 51956 3424
rect 52492 3464 52532 3473
rect 50091 3296 50133 3305
rect 50091 3256 50092 3296
rect 50132 3256 50133 3296
rect 50091 3247 50133 3256
rect 51723 3296 51765 3305
rect 51723 3256 51724 3296
rect 51764 3256 51765 3296
rect 51723 3247 51765 3256
rect 52300 3296 52340 3305
rect 52492 3296 52532 3424
rect 52683 3464 52725 3473
rect 52683 3424 52684 3464
rect 52724 3424 52725 3464
rect 52683 3415 52725 3424
rect 52684 3330 52724 3415
rect 52340 3256 52532 3296
rect 52587 3296 52629 3305
rect 52587 3256 52588 3296
rect 52628 3256 52629 3296
rect 52300 3247 52340 3256
rect 52587 3247 52629 3256
rect 52588 3162 52628 3247
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 3244 2575 3284 2584
rect 3339 2624 3381 2633
rect 3339 2584 3340 2624
rect 3380 2584 3381 2624
rect 3339 2575 3381 2584
rect 6027 2624 6069 2633
rect 6027 2584 6028 2624
rect 6068 2584 6069 2624
rect 6027 2575 6069 2584
rect 3052 2490 3092 2575
rect 3340 2490 3380 2575
rect 53164 2549 53204 5020
rect 53259 5011 53301 5020
rect 53260 4992 53300 5011
rect 53452 4985 53492 7120
rect 53548 7160 53588 7169
rect 53548 6656 53588 7120
rect 53836 6656 53876 6665
rect 53548 6616 53836 6656
rect 53836 6607 53876 6616
rect 53932 6404 53972 8623
rect 53740 6364 53972 6404
rect 54028 8000 54068 8632
rect 54028 6488 54068 7960
rect 54124 8084 54164 8093
rect 54124 7832 54164 8044
rect 54220 8009 54260 8094
rect 54219 8000 54261 8009
rect 54219 7960 54220 8000
rect 54260 7960 54261 8000
rect 54219 7951 54261 7960
rect 54316 8000 54356 9220
rect 54412 8849 54452 9472
rect 54507 9512 54549 9521
rect 54507 9472 54508 9512
rect 54548 9472 54549 9512
rect 54507 9463 54549 9472
rect 54411 8840 54453 8849
rect 54411 8800 54412 8840
rect 54452 8800 54453 8840
rect 54411 8791 54453 8800
rect 54316 7951 54356 7960
rect 54412 8588 54452 8597
rect 54412 7832 54452 8548
rect 54124 7792 54452 7832
rect 54508 7328 54548 9463
rect 54892 9344 54932 9353
rect 54796 8672 54836 8681
rect 54892 8672 54932 9304
rect 54836 8632 54932 8672
rect 54796 8623 54836 8632
rect 55084 8597 55124 10984
rect 56428 11024 56468 11033
rect 56428 10445 56468 10984
rect 56812 11024 56852 11404
rect 56812 10975 56852 10984
rect 56427 10436 56469 10445
rect 56427 10396 56428 10436
rect 56468 10396 56469 10436
rect 56427 10387 56469 10396
rect 56428 9344 56468 9353
rect 55660 8672 55700 8683
rect 55660 8597 55700 8632
rect 55083 8588 55125 8597
rect 55083 8548 55084 8588
rect 55124 8548 55125 8588
rect 55083 8539 55125 8548
rect 55659 8588 55701 8597
rect 55659 8548 55660 8588
rect 55700 8548 55701 8588
rect 55659 8539 55701 8548
rect 55947 8588 55989 8597
rect 55947 8548 55948 8588
rect 55988 8548 55989 8588
rect 55947 8539 55989 8548
rect 55179 8420 55221 8429
rect 55179 8380 55180 8420
rect 55220 8380 55221 8420
rect 55179 8371 55221 8380
rect 55084 7328 55124 7337
rect 54316 7288 54644 7328
rect 54316 7160 54356 7288
rect 54316 7111 54356 7120
rect 54508 7160 54548 7169
rect 54412 7076 54452 7085
rect 54412 6656 54452 7036
rect 54316 6616 54452 6656
rect 54219 6572 54261 6581
rect 54219 6532 54220 6572
rect 54260 6532 54261 6572
rect 54219 6523 54261 6532
rect 54124 6488 54164 6497
rect 54028 6448 54124 6488
rect 53547 5732 53589 5741
rect 53547 5692 53548 5732
rect 53588 5692 53589 5732
rect 53547 5683 53589 5692
rect 53451 4976 53493 4985
rect 53451 4936 53452 4976
rect 53492 4936 53493 4976
rect 53451 4927 53493 4936
rect 53548 4397 53588 5683
rect 53740 5648 53780 6364
rect 53836 6236 53876 6245
rect 53876 6196 53972 6236
rect 53836 6187 53876 6196
rect 53932 5657 53972 6196
rect 53836 5648 53876 5657
rect 53740 5608 53836 5648
rect 53547 4388 53589 4397
rect 53547 4348 53548 4388
rect 53588 4348 53589 4388
rect 53547 4339 53589 4348
rect 53548 4136 53588 4339
rect 53548 4087 53588 4096
rect 53836 3893 53876 5608
rect 53931 5648 53973 5657
rect 53931 5608 53932 5648
rect 53972 5608 53973 5648
rect 53931 5599 53973 5608
rect 54028 4817 54068 6448
rect 54124 6439 54164 6448
rect 54220 6438 54260 6523
rect 54316 6488 54356 6616
rect 54124 5648 54164 5657
rect 54124 5489 54164 5608
rect 54219 5648 54261 5657
rect 54219 5608 54220 5648
rect 54260 5608 54261 5648
rect 54219 5599 54261 5608
rect 54220 5514 54260 5599
rect 54316 5573 54356 6448
rect 54411 6488 54453 6497
rect 54411 6448 54412 6488
rect 54452 6448 54453 6488
rect 54411 6439 54453 6448
rect 54412 6354 54452 6439
rect 54508 5900 54548 7120
rect 54604 6992 54644 7288
rect 54699 7244 54741 7253
rect 54699 7204 54700 7244
rect 54740 7204 54741 7244
rect 54699 7195 54741 7204
rect 54700 7110 54740 7195
rect 54892 6992 54932 7001
rect 54604 6952 54740 6992
rect 54603 6572 54645 6581
rect 54603 6532 54604 6572
rect 54644 6532 54645 6572
rect 54603 6523 54645 6532
rect 54604 6438 54644 6523
rect 54700 6320 54740 6952
rect 54795 6488 54837 6497
rect 54795 6448 54796 6488
rect 54836 6448 54837 6488
rect 54795 6439 54837 6448
rect 54508 5851 54548 5860
rect 54604 6280 54740 6320
rect 54604 5732 54644 6280
rect 54508 5692 54644 5732
rect 54796 5732 54836 6439
rect 54315 5564 54357 5573
rect 54315 5524 54316 5564
rect 54356 5524 54357 5564
rect 54315 5515 54357 5524
rect 54123 5480 54165 5489
rect 54123 5440 54124 5480
rect 54164 5440 54165 5480
rect 54123 5431 54165 5440
rect 54027 4808 54069 4817
rect 54027 4768 54028 4808
rect 54068 4768 54069 4808
rect 54027 4759 54069 4768
rect 53835 3884 53877 3893
rect 53835 3844 53836 3884
rect 53876 3844 53877 3884
rect 53835 3835 53877 3844
rect 53836 3557 53876 3835
rect 53835 3548 53877 3557
rect 53835 3508 53836 3548
rect 53876 3508 53877 3548
rect 53835 3499 53877 3508
rect 54508 3473 54548 5692
rect 54796 5683 54836 5692
rect 54699 5648 54741 5657
rect 54699 5608 54700 5648
rect 54740 5608 54741 5648
rect 54699 5599 54741 5608
rect 54892 5648 54932 6952
rect 54988 6488 55028 6497
rect 55084 6488 55124 7288
rect 55028 6448 55124 6488
rect 54988 6439 55028 6448
rect 54700 5514 54740 5599
rect 54892 5573 54932 5608
rect 54891 5564 54933 5573
rect 54891 5524 54892 5564
rect 54932 5524 54933 5564
rect 54891 5515 54933 5524
rect 54891 4388 54933 4397
rect 54891 4348 54892 4388
rect 54932 4348 54933 4388
rect 54891 4339 54933 4348
rect 54699 4304 54741 4313
rect 54699 4264 54700 4304
rect 54740 4264 54741 4304
rect 54699 4255 54741 4264
rect 54700 4170 54740 4255
rect 54603 4052 54645 4061
rect 54603 4012 54604 4052
rect 54644 4012 54645 4052
rect 54603 4003 54645 4012
rect 54604 3800 54644 4003
rect 54604 3760 54740 3800
rect 54507 3464 54549 3473
rect 54507 3424 54508 3464
rect 54548 3424 54549 3464
rect 54507 3415 54549 3424
rect 53740 3212 53780 3221
rect 53740 2801 53780 3172
rect 53739 2792 53781 2801
rect 53739 2752 53740 2792
rect 53780 2752 53781 2792
rect 53739 2743 53781 2752
rect 53932 2792 53972 2801
rect 53163 2540 53205 2549
rect 53163 2500 53164 2540
rect 53204 2500 53205 2540
rect 53163 2491 53205 2500
rect 1036 2456 1076 2465
rect 1036 2297 1076 2416
rect 1035 2288 1077 2297
rect 1035 2248 1036 2288
rect 1076 2248 1077 2288
rect 1035 2239 1077 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 53452 1952 53492 1961
rect 53452 1793 53492 1912
rect 53836 1952 53876 1961
rect 53932 1952 53972 2752
rect 53876 1912 53972 1952
rect 54700 1952 54740 3760
rect 54892 3464 54932 4339
rect 55180 4313 55220 8371
rect 55948 8084 55988 8539
rect 55948 8035 55988 8044
rect 56332 8000 56372 8009
rect 56428 8000 56468 9304
rect 56811 9008 56853 9017
rect 56811 8968 56812 9008
rect 56852 8968 56853 9008
rect 56811 8959 56853 8968
rect 56812 8924 56852 8959
rect 56812 8873 56852 8884
rect 56372 7960 56468 8000
rect 56332 7951 56372 7960
rect 56812 7076 56852 7085
rect 55852 6488 55892 6497
rect 55852 5741 55892 6448
rect 56812 6329 56852 7036
rect 57004 6656 57044 15259
rect 57195 14888 57237 14897
rect 57195 14848 57196 14888
rect 57236 14848 57237 14888
rect 57195 14839 57237 14848
rect 57100 14720 57140 14729
rect 57100 13721 57140 14680
rect 57196 14720 57236 14839
rect 57196 14671 57236 14680
rect 57099 13712 57141 13721
rect 57099 13672 57100 13712
rect 57140 13672 57141 13712
rect 57099 13663 57141 13672
rect 57292 12980 57332 16015
rect 57484 15560 57524 16360
rect 57580 16351 57620 16360
rect 57964 16232 58004 17107
rect 58055 17072 58095 17472
rect 58345 17249 58385 17472
rect 58344 17240 58386 17249
rect 58252 17200 58345 17240
rect 58385 17200 58386 17240
rect 58055 17032 58100 17072
rect 58060 16484 58100 17032
rect 58060 16435 58100 16444
rect 57964 16183 58004 16192
rect 58252 16232 58292 17200
rect 58344 17191 58386 17200
rect 58455 17072 58495 17472
rect 58745 17156 58785 17472
rect 58348 17032 58495 17072
rect 58540 17116 58785 17156
rect 58348 16484 58388 17032
rect 58348 16435 58388 16444
rect 58540 16241 58580 17116
rect 58855 17072 58895 17472
rect 59145 17156 59185 17472
rect 58636 17032 58895 17072
rect 59116 17116 59185 17156
rect 58636 16484 58676 17032
rect 58636 16435 58676 16444
rect 58252 16183 58292 16192
rect 58539 16232 58581 16241
rect 58539 16192 58540 16232
rect 58580 16192 58581 16232
rect 58539 16183 58581 16192
rect 58924 16232 58964 16241
rect 59116 16232 59156 17116
rect 59255 17072 59295 17472
rect 59545 17156 59585 17472
rect 58964 16192 59156 16232
rect 59212 17032 59295 17072
rect 59500 17116 59585 17156
rect 58540 16098 58580 16183
rect 58924 15821 58964 16192
rect 59020 16064 59060 16073
rect 59212 16064 59252 17032
rect 59060 16024 59252 16064
rect 59308 16232 59348 16241
rect 59500 16232 59540 17116
rect 59655 17072 59695 17472
rect 59945 17156 59985 17472
rect 59348 16192 59540 16232
rect 59596 17032 59695 17072
rect 59884 17116 59985 17156
rect 59020 16015 59060 16024
rect 58923 15812 58965 15821
rect 58923 15772 58924 15812
rect 58964 15772 58965 15812
rect 58923 15763 58965 15772
rect 57484 15511 57524 15520
rect 58348 15560 58388 15569
rect 57483 14888 57525 14897
rect 57483 14848 57484 14888
rect 57524 14848 57525 14888
rect 57483 14839 57525 14848
rect 57484 14754 57524 14839
rect 57388 14720 57428 14729
rect 57388 13469 57428 14680
rect 57579 14720 57621 14729
rect 57579 14680 57580 14720
rect 57620 14680 57621 14720
rect 57579 14671 57621 14680
rect 57580 14586 57620 14671
rect 57675 14636 57717 14645
rect 57675 14596 57676 14636
rect 57716 14596 57717 14636
rect 57675 14587 57717 14596
rect 57387 13460 57429 13469
rect 57387 13420 57388 13460
rect 57428 13420 57429 13460
rect 57387 13411 57429 13420
rect 57676 13208 57716 14587
rect 58348 14477 58388 15520
rect 58636 14888 58676 14897
rect 58540 14848 58636 14888
rect 58347 14468 58389 14477
rect 58347 14428 58348 14468
rect 58388 14428 58389 14468
rect 58347 14419 58389 14428
rect 57963 14300 58005 14309
rect 57963 14260 57964 14300
rect 58004 14260 58005 14300
rect 57963 14251 58005 14260
rect 57771 14048 57813 14057
rect 57771 14008 57772 14048
rect 57812 14008 57813 14048
rect 57771 13999 57813 14008
rect 57964 14048 58004 14251
rect 58156 14048 58196 14057
rect 58540 14048 58580 14848
rect 58636 14839 58676 14848
rect 58827 14552 58869 14561
rect 58827 14512 58828 14552
rect 58868 14512 58869 14552
rect 58827 14503 58869 14512
rect 58004 14008 58100 14048
rect 57964 13999 58004 14008
rect 57772 13914 57812 13999
rect 57867 13796 57909 13805
rect 57867 13756 57868 13796
rect 57908 13756 57909 13796
rect 57867 13747 57909 13756
rect 57868 13662 57908 13747
rect 57963 13544 58005 13553
rect 57963 13504 57964 13544
rect 58004 13504 58005 13544
rect 57963 13495 58005 13504
rect 57868 13208 57908 13217
rect 57676 13168 57868 13208
rect 57868 13159 57908 13168
rect 57675 13040 57717 13049
rect 57675 13000 57676 13040
rect 57716 13000 57717 13040
rect 57675 12991 57717 13000
rect 57867 13040 57909 13049
rect 57867 13000 57868 13040
rect 57908 13000 57909 13040
rect 57867 12991 57909 13000
rect 57196 12940 57332 12980
rect 57196 9185 57236 12940
rect 57291 12704 57333 12713
rect 57291 12664 57292 12704
rect 57332 12664 57333 12704
rect 57291 12655 57333 12664
rect 57292 12570 57332 12655
rect 57579 12536 57621 12545
rect 57579 12496 57580 12536
rect 57620 12496 57621 12536
rect 57579 12487 57621 12496
rect 57483 12032 57525 12041
rect 57483 11992 57484 12032
rect 57524 11992 57525 12032
rect 57483 11983 57525 11992
rect 57292 11864 57332 11873
rect 57292 11621 57332 11824
rect 57484 11780 57524 11983
rect 57484 11731 57524 11740
rect 57291 11612 57333 11621
rect 57291 11572 57292 11612
rect 57332 11572 57333 11612
rect 57291 11563 57333 11572
rect 57292 9428 57332 11563
rect 57580 11024 57620 12487
rect 57676 11696 57716 12991
rect 57868 12452 57908 12991
rect 57868 12403 57908 12412
rect 57964 12284 58004 13495
rect 58060 13208 58100 14008
rect 58196 14008 58484 14048
rect 58156 13999 58196 14008
rect 58347 13880 58389 13889
rect 58347 13840 58348 13880
rect 58388 13840 58389 13880
rect 58347 13831 58389 13840
rect 58156 13208 58196 13217
rect 58060 13168 58156 13208
rect 58156 13159 58196 13168
rect 58252 13124 58292 13133
rect 58252 12713 58292 13084
rect 58251 12704 58293 12713
rect 58156 12664 58252 12704
rect 58292 12664 58293 12704
rect 57676 11647 57716 11656
rect 57868 12244 58004 12284
rect 58059 12284 58101 12293
rect 58059 12244 58060 12284
rect 58100 12244 58101 12284
rect 57868 11696 57908 12244
rect 58059 12235 58101 12244
rect 58060 12150 58100 12235
rect 58156 11789 58196 12664
rect 58251 12655 58293 12664
rect 58252 12536 58292 12545
rect 58348 12536 58388 13831
rect 58444 13544 58484 14008
rect 58540 13999 58580 14008
rect 58444 13504 58772 13544
rect 58732 13460 58772 13504
rect 58732 13411 58772 13420
rect 58540 13376 58580 13385
rect 58292 12496 58388 12536
rect 58444 13336 58540 13376
rect 58444 12536 58484 13336
rect 58540 13327 58580 13336
rect 58539 13208 58581 13217
rect 58539 13168 58540 13208
rect 58580 13168 58581 13208
rect 58539 13159 58581 13168
rect 58732 13208 58772 13217
rect 58828 13208 58868 14503
rect 59019 13796 59061 13805
rect 59019 13756 59020 13796
rect 59060 13756 59061 13796
rect 59019 13747 59061 13756
rect 58772 13168 58868 13208
rect 58923 13208 58965 13217
rect 58923 13168 58924 13208
rect 58964 13168 58965 13208
rect 58732 13159 58772 13168
rect 58923 13159 58965 13168
rect 59020 13208 59060 13747
rect 59020 13159 59060 13168
rect 58252 12487 58292 12496
rect 58444 12487 58484 12496
rect 58348 12368 58388 12377
rect 58540 12368 58580 13159
rect 58924 13074 58964 13159
rect 59308 12797 59348 16192
rect 59596 16148 59636 17032
rect 59404 16108 59636 16148
rect 59692 16232 59732 16241
rect 59884 16232 59924 17116
rect 60055 17072 60095 17472
rect 60345 17072 60385 17472
rect 59732 16192 59924 16232
rect 59980 17032 60095 17072
rect 60268 17032 60385 17072
rect 59404 16064 59444 16108
rect 59404 16015 59444 16024
rect 59499 15980 59541 15989
rect 59499 15940 59500 15980
rect 59540 15940 59541 15980
rect 59499 15931 59541 15940
rect 59500 15728 59540 15931
rect 59500 15679 59540 15688
rect 59500 15308 59540 15317
rect 59500 14729 59540 15268
rect 59499 14720 59541 14729
rect 59499 14680 59500 14720
rect 59540 14680 59541 14720
rect 59499 14671 59541 14680
rect 59499 14552 59541 14561
rect 59499 14512 59500 14552
rect 59540 14512 59541 14552
rect 59499 14503 59541 14512
rect 59403 14384 59445 14393
rect 59403 14344 59404 14384
rect 59444 14344 59445 14384
rect 59403 14335 59445 14344
rect 59404 14048 59444 14335
rect 59404 13999 59444 14008
rect 59307 12788 59349 12797
rect 59307 12748 59308 12788
rect 59348 12748 59349 12788
rect 59307 12739 59349 12748
rect 59307 12620 59349 12629
rect 59307 12580 59308 12620
rect 59348 12580 59349 12620
rect 59307 12571 59349 12580
rect 59019 12536 59061 12545
rect 59019 12496 59020 12536
rect 59060 12496 59061 12536
rect 59019 12487 59061 12496
rect 59308 12536 59348 12571
rect 58388 12328 58580 12368
rect 58348 12319 58388 12328
rect 58251 12284 58293 12293
rect 58251 12244 58252 12284
rect 58292 12244 58293 12284
rect 58251 12235 58293 12244
rect 58252 11948 58292 12235
rect 59020 12125 59060 12487
rect 59115 12284 59157 12293
rect 59115 12244 59116 12284
rect 59156 12244 59157 12284
rect 59115 12235 59157 12244
rect 59019 12116 59061 12125
rect 59019 12076 59020 12116
rect 59060 12076 59061 12116
rect 59019 12067 59061 12076
rect 58252 11908 58676 11948
rect 57963 11780 58005 11789
rect 57963 11740 57964 11780
rect 58004 11740 58005 11780
rect 57963 11731 58005 11740
rect 58155 11780 58197 11789
rect 58155 11740 58156 11780
rect 58196 11740 58197 11780
rect 58155 11731 58197 11740
rect 57868 11647 57908 11656
rect 57964 11696 58004 11731
rect 57964 11645 58004 11656
rect 58252 11696 58292 11908
rect 58348 11789 58388 11820
rect 58347 11780 58389 11789
rect 58347 11740 58348 11780
rect 58388 11740 58389 11780
rect 58347 11731 58389 11740
rect 58252 11647 58292 11656
rect 58348 11696 58388 11731
rect 58348 11621 58388 11656
rect 58444 11696 58484 11705
rect 58347 11612 58389 11621
rect 58347 11572 58348 11612
rect 58388 11572 58389 11612
rect 58347 11563 58389 11572
rect 57772 11528 57812 11537
rect 57676 11024 57716 11033
rect 57580 10984 57676 11024
rect 57676 10975 57716 10984
rect 57579 10352 57621 10361
rect 57579 10312 57580 10352
rect 57620 10312 57621 10352
rect 57579 10303 57621 10312
rect 57387 10268 57429 10277
rect 57387 10228 57388 10268
rect 57428 10228 57429 10268
rect 57387 10219 57429 10228
rect 57388 10134 57428 10219
rect 57580 10218 57620 10303
rect 57772 10184 57812 11488
rect 58156 11528 58196 11537
rect 58059 10436 58101 10445
rect 58059 10396 58060 10436
rect 58100 10396 58101 10436
rect 58059 10387 58101 10396
rect 58060 10302 58100 10387
rect 57772 10135 57812 10144
rect 57867 10184 57909 10193
rect 57867 10144 57868 10184
rect 57908 10144 57909 10184
rect 57867 10135 57909 10144
rect 58060 10184 58100 10193
rect 58156 10184 58196 11488
rect 58444 11201 58484 11656
rect 58443 11192 58485 11201
rect 58443 11152 58444 11192
rect 58484 11152 58580 11192
rect 58443 11143 58485 11152
rect 58251 10352 58293 10361
rect 58251 10312 58252 10352
rect 58292 10312 58293 10352
rect 58251 10303 58293 10312
rect 58100 10144 58196 10184
rect 58252 10184 58292 10303
rect 58060 10135 58100 10144
rect 57868 10050 57908 10135
rect 58059 10016 58101 10025
rect 58059 9976 58060 10016
rect 58100 9976 58101 10016
rect 58059 9967 58101 9976
rect 57772 9512 57812 9521
rect 57676 9472 57772 9512
rect 57388 9428 57428 9437
rect 57292 9388 57388 9428
rect 57388 9379 57428 9388
rect 57580 9260 57620 9269
rect 57195 9176 57237 9185
rect 57195 9136 57196 9176
rect 57236 9136 57237 9176
rect 57195 9127 57237 9136
rect 57580 8336 57620 9220
rect 57676 8672 57716 9472
rect 57772 9463 57812 9472
rect 57964 9512 58004 9521
rect 57772 9260 57812 9269
rect 57772 8849 57812 9220
rect 57964 8849 58004 9472
rect 58060 9512 58100 9967
rect 58252 9932 58292 10144
rect 58444 10184 58484 10193
rect 58347 10016 58389 10025
rect 58347 9976 58348 10016
rect 58388 9976 58389 10016
rect 58347 9967 58389 9976
rect 58060 9463 58100 9472
rect 58156 9892 58292 9932
rect 58059 9092 58101 9101
rect 58059 9052 58060 9092
rect 58100 9052 58101 9092
rect 58059 9043 58101 9052
rect 57771 8840 57813 8849
rect 57771 8800 57772 8840
rect 57812 8800 57813 8840
rect 57771 8791 57813 8800
rect 57963 8840 58005 8849
rect 57963 8800 57964 8840
rect 58004 8800 58005 8840
rect 57963 8791 58005 8800
rect 57772 8672 57812 8681
rect 57676 8632 57772 8672
rect 57772 8623 57812 8632
rect 57868 8672 57908 8681
rect 57868 8513 57908 8632
rect 57964 8672 58004 8681
rect 57867 8504 57909 8513
rect 57867 8464 57868 8504
rect 57908 8464 57909 8504
rect 57867 8455 57909 8464
rect 57964 8336 58004 8632
rect 58060 8672 58100 9043
rect 58060 8623 58100 8632
rect 57580 8296 58004 8336
rect 57196 8000 57236 8009
rect 57236 7960 57428 8000
rect 57196 7951 57236 7960
rect 57004 6607 57044 6616
rect 57196 7160 57236 7169
rect 56811 6320 56853 6329
rect 56811 6280 56812 6320
rect 56852 6280 56853 6320
rect 57196 6320 57236 7120
rect 57292 6320 57332 6329
rect 57196 6280 57292 6320
rect 56811 6271 56853 6280
rect 57292 6271 57332 6280
rect 57004 6236 57044 6245
rect 56620 5816 56660 5825
rect 55851 5732 55893 5741
rect 55851 5692 55852 5732
rect 55892 5692 55893 5732
rect 55851 5683 55893 5692
rect 56236 5648 56276 5659
rect 56236 5573 56276 5608
rect 56428 5648 56468 5657
rect 56235 5564 56277 5573
rect 56235 5524 56236 5564
rect 56276 5524 56277 5564
rect 56235 5515 56277 5524
rect 56332 5564 56372 5573
rect 55756 5144 55796 5153
rect 55796 5104 56084 5144
rect 55756 5095 55796 5104
rect 56044 5060 56084 5104
rect 56140 5060 56180 5069
rect 56044 5020 56140 5060
rect 56140 5011 56180 5020
rect 55660 4976 55700 4985
rect 55660 4817 55700 4936
rect 55852 4976 55892 4985
rect 55659 4808 55701 4817
rect 55659 4768 55660 4808
rect 55700 4768 55701 4808
rect 55659 4759 55701 4768
rect 55852 4397 55892 4936
rect 55947 4976 55989 4985
rect 55947 4936 55948 4976
rect 55988 4936 55989 4976
rect 55947 4927 55989 4936
rect 55948 4842 55988 4927
rect 55851 4388 55893 4397
rect 56236 4388 56276 5515
rect 56332 4985 56372 5524
rect 56331 4976 56373 4985
rect 56331 4936 56332 4976
rect 56372 4936 56373 4976
rect 56331 4927 56373 4936
rect 56331 4808 56373 4817
rect 56331 4768 56332 4808
rect 56372 4768 56373 4808
rect 56331 4759 56373 4768
rect 55851 4348 55852 4388
rect 55892 4348 55893 4388
rect 55851 4339 55893 4348
rect 56044 4348 56276 4388
rect 55084 4304 55124 4313
rect 55084 3809 55124 4264
rect 55179 4304 55221 4313
rect 55179 4264 55180 4304
rect 55220 4264 55221 4304
rect 55179 4255 55221 4264
rect 55659 4220 55701 4229
rect 55659 4180 55660 4220
rect 55700 4180 55701 4220
rect 55659 4171 55701 4180
rect 55563 4136 55605 4145
rect 55563 4096 55564 4136
rect 55604 4096 55605 4136
rect 55563 4087 55605 4096
rect 55660 4136 55700 4171
rect 55564 4002 55604 4087
rect 55083 3800 55125 3809
rect 55083 3760 55084 3800
rect 55124 3760 55125 3800
rect 55083 3751 55125 3760
rect 55660 3548 55700 4096
rect 55756 4136 55796 4145
rect 55756 3977 55796 4096
rect 55852 4136 55892 4145
rect 55852 4052 55892 4096
rect 55852 4012 55979 4052
rect 55939 3977 55979 4012
rect 55755 3968 55797 3977
rect 55939 3968 55989 3977
rect 55755 3928 55756 3968
rect 55796 3928 55892 3968
rect 55939 3928 55948 3968
rect 55988 3928 55989 3968
rect 55755 3919 55797 3928
rect 55755 3800 55797 3809
rect 55755 3760 55756 3800
rect 55796 3760 55797 3800
rect 55755 3751 55797 3760
rect 54892 3415 54932 3424
rect 55564 3508 55700 3548
rect 55467 2204 55509 2213
rect 55467 2164 55468 2204
rect 55508 2164 55509 2204
rect 55467 2155 55509 2164
rect 53836 1903 53876 1912
rect 54700 1903 54740 1912
rect 53451 1784 53493 1793
rect 53451 1744 53452 1784
rect 53492 1744 53493 1784
rect 53451 1735 53493 1744
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 55468 1112 55508 2155
rect 55468 1063 55508 1072
rect 55564 1112 55604 3508
rect 55756 3464 55796 3751
rect 55756 3415 55796 3424
rect 55852 3296 55892 3928
rect 55947 3919 55989 3928
rect 55564 1063 55604 1072
rect 55660 3256 55892 3296
rect 55660 1112 55700 3256
rect 55948 3212 55988 3919
rect 55756 3172 55988 3212
rect 55756 2801 55796 3172
rect 56044 2900 56084 4348
rect 56140 4136 56180 4145
rect 56140 3893 56180 4096
rect 56139 3884 56181 3893
rect 56139 3844 56140 3884
rect 56180 3844 56181 3884
rect 56139 3835 56181 3844
rect 56140 3716 56180 3835
rect 56140 3676 56276 3716
rect 56139 3548 56181 3557
rect 56139 3508 56140 3548
rect 56180 3508 56181 3548
rect 56139 3499 56181 3508
rect 56140 3414 56180 3499
rect 56236 3296 56276 3676
rect 55852 2860 56084 2900
rect 56140 3256 56276 3296
rect 55755 2792 55797 2801
rect 55755 2752 55756 2792
rect 55796 2752 55797 2792
rect 55755 2743 55797 2752
rect 55756 2624 55796 2743
rect 55852 2717 55892 2860
rect 55851 2708 55893 2717
rect 55851 2668 55852 2708
rect 55892 2668 55893 2708
rect 55851 2659 55893 2668
rect 55756 2575 55796 2584
rect 55852 2624 55892 2659
rect 55852 2574 55892 2584
rect 56044 2582 56084 2591
rect 56043 2542 56044 2549
rect 56084 2542 56085 2549
rect 56043 2540 56085 2542
rect 56043 2500 56044 2540
rect 56084 2500 56085 2540
rect 56043 2491 56085 2500
rect 55948 2456 55988 2465
rect 56044 2447 56084 2491
rect 55851 2120 55893 2129
rect 55851 2080 55852 2120
rect 55892 2080 55893 2120
rect 55851 2071 55893 2080
rect 55852 1986 55892 2071
rect 55948 1961 55988 2416
rect 56043 2204 56085 2213
rect 56043 2164 56044 2204
rect 56084 2164 56085 2204
rect 56043 2155 56085 2164
rect 55947 1952 55989 1961
rect 55947 1912 55948 1952
rect 55988 1912 55989 1952
rect 55947 1903 55989 1912
rect 56044 1952 56084 2155
rect 56044 1903 56084 1912
rect 55947 1784 55989 1793
rect 56044 1784 56084 1793
rect 55947 1744 55948 1784
rect 55988 1744 56044 1784
rect 55947 1735 55989 1744
rect 56044 1735 56084 1744
rect 55755 1196 55797 1205
rect 55755 1156 55756 1196
rect 55796 1156 55797 1196
rect 55755 1147 55797 1156
rect 55660 1063 55700 1072
rect 55756 1112 55796 1147
rect 55756 1061 55796 1072
rect 56140 1112 56180 3256
rect 56235 2792 56277 2801
rect 56235 2752 56236 2792
rect 56276 2752 56277 2792
rect 56235 2743 56277 2752
rect 56236 1952 56276 2743
rect 56332 2624 56372 4759
rect 56428 4733 56468 5608
rect 56524 4976 56564 4985
rect 56620 4976 56660 5776
rect 57004 5657 57044 6196
rect 57388 5741 57428 7960
rect 57771 6824 57813 6833
rect 57771 6784 57772 6824
rect 57812 6784 57813 6824
rect 57771 6775 57813 6784
rect 57387 5732 57429 5741
rect 57387 5692 57388 5732
rect 57428 5692 57429 5732
rect 57387 5683 57429 5692
rect 57003 5648 57045 5657
rect 57003 5608 57004 5648
rect 57044 5608 57045 5648
rect 57003 5599 57045 5608
rect 56564 4936 56660 4976
rect 57388 4976 57428 5683
rect 56524 4927 56564 4936
rect 57388 4927 57428 4936
rect 56427 4724 56469 4733
rect 56427 4684 56428 4724
rect 56468 4684 56469 4724
rect 56427 4675 56469 4684
rect 56428 4136 56468 4675
rect 56715 4388 56757 4397
rect 56715 4348 56716 4388
rect 56756 4348 56757 4388
rect 56715 4339 56757 4348
rect 57195 4388 57237 4397
rect 57195 4348 57196 4388
rect 57236 4348 57237 4388
rect 57772 4388 57812 6775
rect 57868 6413 57908 8296
rect 58156 8009 58196 9892
rect 58348 9882 58388 9967
rect 58348 9512 58388 9521
rect 58348 9185 58388 9472
rect 58347 9176 58389 9185
rect 58347 9136 58348 9176
rect 58388 9136 58389 9176
rect 58347 9127 58389 9136
rect 58251 9092 58293 9101
rect 58251 9052 58252 9092
rect 58292 9052 58293 9092
rect 58251 9043 58293 9052
rect 58252 8924 58292 9043
rect 58252 8884 58388 8924
rect 58251 8756 58293 8765
rect 58251 8716 58252 8756
rect 58292 8716 58293 8756
rect 58251 8707 58293 8716
rect 58252 8622 58292 8707
rect 58348 8168 58388 8884
rect 58444 8672 58484 10144
rect 58540 10184 58580 11152
rect 58540 10135 58580 10144
rect 58636 10016 58676 11908
rect 58827 11696 58869 11705
rect 58732 11656 58828 11696
rect 58868 11656 58869 11696
rect 58732 10940 58772 11656
rect 58827 11647 58869 11656
rect 59020 11696 59060 11705
rect 58828 11562 58868 11647
rect 58923 11612 58965 11621
rect 58923 11572 58924 11612
rect 58964 11572 58965 11612
rect 58923 11563 58965 11572
rect 58924 11478 58964 11563
rect 58827 11192 58869 11201
rect 58827 11152 58828 11192
rect 58868 11152 58869 11192
rect 58827 11143 58869 11152
rect 58828 11058 58868 11143
rect 59020 10940 59060 11656
rect 59116 11696 59156 12235
rect 59308 11948 59348 12496
rect 59500 12536 59540 14503
rect 59692 12545 59732 16192
rect 59788 16064 59828 16073
rect 59980 16064 60020 17032
rect 60268 16988 60308 17032
rect 60455 16988 60495 17472
rect 60745 17156 60785 17472
rect 59828 16024 60020 16064
rect 60076 16948 60308 16988
rect 60364 16948 60495 16988
rect 60556 17116 60785 17156
rect 60076 16232 60116 16948
rect 60172 16484 60212 16493
rect 60364 16484 60404 16948
rect 60212 16444 60404 16484
rect 60172 16435 60212 16444
rect 59788 16015 59828 16024
rect 59691 12536 59733 12545
rect 59540 12496 59636 12536
rect 59500 12487 59540 12496
rect 59403 12284 59445 12293
rect 59403 12244 59404 12284
rect 59444 12244 59445 12284
rect 59403 12235 59445 12244
rect 59404 12150 59444 12235
rect 59308 11908 59444 11948
rect 59116 11647 59156 11656
rect 59307 11612 59349 11621
rect 59307 11572 59308 11612
rect 59348 11572 59349 11612
rect 59307 11563 59349 11572
rect 59308 11478 59348 11563
rect 59307 11192 59349 11201
rect 59307 11152 59308 11192
rect 59348 11152 59349 11192
rect 59307 11143 59349 11152
rect 59308 11108 59348 11143
rect 59308 11057 59348 11068
rect 59404 11024 59444 11908
rect 59499 11528 59541 11537
rect 59499 11488 59500 11528
rect 59540 11488 59541 11528
rect 59596 11528 59636 12496
rect 59691 12496 59692 12536
rect 59732 12496 59733 12536
rect 59691 12487 59733 12496
rect 59788 12368 59828 12377
rect 59692 12328 59788 12368
rect 59692 11696 59732 12328
rect 59788 12319 59828 12328
rect 59692 11647 59732 11656
rect 59596 11488 59828 11528
rect 59499 11479 59541 11488
rect 59404 10975 59444 10984
rect 58732 10900 58868 10940
rect 59020 10900 59156 10940
rect 58732 10352 58772 10363
rect 58732 10277 58772 10312
rect 58731 10268 58773 10277
rect 58731 10228 58732 10268
rect 58772 10228 58773 10268
rect 58731 10219 58773 10228
rect 58540 9976 58676 10016
rect 58540 8849 58580 9976
rect 58636 9512 58676 9521
rect 58636 9353 58676 9472
rect 58732 9512 58772 9521
rect 58635 9344 58677 9353
rect 58635 9304 58636 9344
rect 58676 9304 58677 9344
rect 58635 9295 58677 9304
rect 58732 9101 58772 9472
rect 58731 9092 58773 9101
rect 58731 9052 58732 9092
rect 58772 9052 58773 9092
rect 58731 9043 58773 9052
rect 58539 8840 58581 8849
rect 58539 8800 58540 8840
rect 58580 8800 58581 8840
rect 58539 8791 58581 8800
rect 58732 8756 58772 8765
rect 58828 8756 58868 10900
rect 59020 10772 59060 10781
rect 58923 10268 58965 10277
rect 58923 10228 58924 10268
rect 58964 10228 58965 10268
rect 58923 10219 58965 10228
rect 58924 10134 58964 10219
rect 59020 10184 59060 10732
rect 59116 10352 59156 10900
rect 59116 10312 59252 10352
rect 59212 10193 59252 10312
rect 59500 10268 59540 11479
rect 59691 11024 59733 11033
rect 59116 10184 59156 10193
rect 59020 10144 59116 10184
rect 59116 10135 59156 10144
rect 59211 10184 59253 10193
rect 59211 10144 59212 10184
rect 59252 10144 59253 10184
rect 59211 10135 59253 10144
rect 59308 10184 59348 10193
rect 59500 10184 59540 10228
rect 59348 10144 59540 10184
rect 59596 10984 59692 11024
rect 59732 10984 59733 11024
rect 59308 10135 59348 10144
rect 59212 10100 59252 10135
rect 59596 10100 59636 10984
rect 59691 10975 59733 10984
rect 59692 10890 59732 10975
rect 59788 10268 59828 11488
rect 60076 10865 60116 16192
rect 60171 16232 60213 16241
rect 60556 16232 60596 17116
rect 60855 17072 60895 17472
rect 61145 17072 61185 17472
rect 60652 17032 60895 17072
rect 61132 17032 61185 17072
rect 61255 17072 61295 17472
rect 61545 17249 61585 17472
rect 61544 17240 61586 17249
rect 61544 17200 61545 17240
rect 61585 17200 61586 17240
rect 61544 17191 61586 17200
rect 61655 17072 61695 17472
rect 61945 17324 61985 17472
rect 61900 17284 61985 17324
rect 61803 17240 61845 17249
rect 61803 17200 61804 17240
rect 61844 17200 61845 17240
rect 61803 17191 61845 17200
rect 61255 17032 61556 17072
rect 61655 17032 61748 17072
rect 60652 16484 60692 17032
rect 60652 16435 60692 16444
rect 60171 16192 60172 16232
rect 60212 16192 60213 16232
rect 60171 16183 60213 16192
rect 60364 16192 60556 16232
rect 60075 10856 60117 10865
rect 60075 10816 60076 10856
rect 60116 10816 60117 10856
rect 60075 10807 60117 10816
rect 60076 10268 60116 10277
rect 59788 10228 60076 10268
rect 60076 10219 60116 10228
rect 59212 10050 59252 10060
rect 59404 10060 59636 10100
rect 59883 10100 59925 10109
rect 59883 10060 59884 10100
rect 59924 10060 59925 10100
rect 59404 9428 59444 10060
rect 59883 10051 59925 10060
rect 59692 10016 59732 10025
rect 59884 10016 59924 10051
rect 59732 9976 59828 10016
rect 59692 9967 59732 9976
rect 59596 9512 59636 9521
rect 59404 9379 59444 9388
rect 59500 9472 59596 9512
rect 59020 9260 59060 9269
rect 59020 8933 59060 9220
rect 59212 9260 59252 9271
rect 59212 9185 59252 9220
rect 59307 9260 59349 9269
rect 59307 9220 59308 9260
rect 59348 9220 59349 9260
rect 59307 9211 59349 9220
rect 59211 9176 59253 9185
rect 59211 9136 59212 9176
rect 59252 9136 59253 9176
rect 59211 9127 59253 9136
rect 59308 9101 59348 9211
rect 59307 9092 59349 9101
rect 59307 9052 59308 9092
rect 59348 9052 59349 9092
rect 59307 9043 59349 9052
rect 59019 8924 59061 8933
rect 59019 8884 59020 8924
rect 59060 8884 59061 8924
rect 59019 8875 59061 8884
rect 58772 8716 58868 8756
rect 58924 8840 58964 8849
rect 59500 8840 59540 9472
rect 59596 9463 59636 9472
rect 59691 8924 59733 8933
rect 58732 8707 58772 8716
rect 58924 8672 58964 8800
rect 59212 8800 59540 8840
rect 59596 8884 59692 8924
rect 59732 8884 59733 8924
rect 59116 8672 59156 8681
rect 58444 8632 58676 8672
rect 58443 8504 58485 8513
rect 58443 8464 58444 8504
rect 58484 8464 58485 8504
rect 58443 8455 58485 8464
rect 58444 8370 58484 8455
rect 58388 8128 58580 8168
rect 58348 8119 58388 8128
rect 58155 8000 58197 8009
rect 58155 7960 58156 8000
rect 58196 7960 58197 8000
rect 58155 7951 58197 7960
rect 58540 8000 58580 8128
rect 58540 7951 58580 7960
rect 58636 8000 58676 8632
rect 58924 8632 59116 8672
rect 58731 8504 58773 8513
rect 58731 8464 58732 8504
rect 58772 8464 58773 8504
rect 58731 8455 58773 8464
rect 58636 7832 58676 7960
rect 58252 7792 58676 7832
rect 58060 7160 58100 7169
rect 57964 7120 58060 7160
rect 57867 6404 57909 6413
rect 57867 6364 57868 6404
rect 57908 6364 57909 6404
rect 57867 6355 57909 6364
rect 57964 5741 58004 7120
rect 58060 7111 58100 7120
rect 58252 6740 58292 7792
rect 58156 6700 58292 6740
rect 58060 6497 58100 6582
rect 58059 6488 58101 6497
rect 58059 6448 58060 6488
rect 58100 6448 58101 6488
rect 58059 6439 58101 6448
rect 58059 6320 58101 6329
rect 58059 6280 58060 6320
rect 58100 6280 58101 6320
rect 58059 6271 58101 6280
rect 58060 6186 58100 6271
rect 57963 5732 58005 5741
rect 57963 5692 57964 5732
rect 58004 5692 58005 5732
rect 57963 5683 58005 5692
rect 58156 5573 58196 6700
rect 58347 6656 58389 6665
rect 58732 6656 58772 8455
rect 58827 8000 58869 8009
rect 58827 7960 58828 8000
rect 58868 7960 58869 8000
rect 58827 7951 58869 7960
rect 58828 7866 58868 7951
rect 58828 7748 58868 7757
rect 58828 6665 58868 7708
rect 58924 7169 58964 8632
rect 59116 8623 59156 8632
rect 59212 8588 59252 8800
rect 59308 8672 59348 8683
rect 59308 8597 59348 8632
rect 59403 8672 59445 8681
rect 59403 8632 59404 8672
rect 59444 8632 59445 8672
rect 59403 8623 59445 8632
rect 59596 8672 59636 8884
rect 59691 8875 59733 8884
rect 59691 8756 59733 8765
rect 59691 8716 59692 8756
rect 59732 8716 59733 8756
rect 59691 8707 59733 8716
rect 59596 8623 59636 8632
rect 59212 8539 59252 8548
rect 59307 8588 59349 8597
rect 59307 8548 59308 8588
rect 59348 8548 59349 8588
rect 59307 8539 59349 8548
rect 59404 8538 59444 8623
rect 59692 8622 59732 8707
rect 59788 8672 59828 9976
rect 59884 9344 59924 9976
rect 59979 10016 60021 10025
rect 59979 9976 59980 10016
rect 60020 9976 60021 10016
rect 59979 9967 60021 9976
rect 59980 9512 60020 9967
rect 59980 9463 60020 9472
rect 60172 9428 60212 16183
rect 60364 10529 60404 16192
rect 60556 16183 60596 16192
rect 61036 16400 61076 16409
rect 60556 15560 60596 15569
rect 60940 15560 60980 15569
rect 61036 15560 61076 16360
rect 61132 16073 61172 17032
rect 61516 16484 61556 17032
rect 61708 16493 61748 17032
rect 61516 16435 61556 16444
rect 61707 16484 61749 16493
rect 61707 16444 61708 16484
rect 61748 16444 61749 16484
rect 61707 16435 61749 16444
rect 61707 16316 61749 16325
rect 61707 16276 61708 16316
rect 61748 16276 61749 16316
rect 61707 16267 61749 16276
rect 61420 16232 61460 16241
rect 61420 16073 61460 16192
rect 61708 16182 61748 16267
rect 61611 16148 61653 16157
rect 61611 16108 61612 16148
rect 61652 16108 61653 16148
rect 61611 16099 61653 16108
rect 61131 16064 61173 16073
rect 61131 16024 61132 16064
rect 61172 16024 61173 16064
rect 61131 16015 61173 16024
rect 61419 16064 61461 16073
rect 61419 16024 61420 16064
rect 61460 16024 61461 16064
rect 61419 16015 61461 16024
rect 60596 15520 60788 15560
rect 60556 15511 60596 15520
rect 60748 14972 60788 15520
rect 60980 15520 61076 15560
rect 60940 15511 60980 15520
rect 61612 15317 61652 16099
rect 61804 15905 61844 17191
rect 61900 16241 61940 17284
rect 62055 17072 62095 17472
rect 62345 17249 62385 17472
rect 62344 17240 62386 17249
rect 62344 17200 62345 17240
rect 62385 17200 62386 17240
rect 62344 17191 62386 17200
rect 62455 17072 62495 17472
rect 62745 17156 62785 17472
rect 62745 17116 62804 17156
rect 62667 17072 62709 17081
rect 62055 17032 62324 17072
rect 62455 17032 62612 17072
rect 62187 16484 62229 16493
rect 62187 16444 62188 16484
rect 62228 16444 62229 16484
rect 62284 16484 62324 17032
rect 62476 16484 62516 16493
rect 62284 16444 62476 16484
rect 62187 16435 62229 16444
rect 62476 16435 62516 16444
rect 62188 16350 62228 16435
rect 61899 16232 61941 16241
rect 61899 16192 61900 16232
rect 61940 16192 61941 16232
rect 61899 16183 61941 16192
rect 62092 16232 62132 16241
rect 61900 16064 61940 16073
rect 61940 16024 62036 16064
rect 61900 16015 61940 16024
rect 61803 15896 61845 15905
rect 61803 15856 61804 15896
rect 61844 15856 61845 15896
rect 61803 15847 61845 15856
rect 61996 15569 62036 16024
rect 62092 15905 62132 16192
rect 62379 16232 62421 16241
rect 62379 16192 62380 16232
rect 62420 16192 62421 16232
rect 62379 16183 62421 16192
rect 62380 16098 62420 16183
rect 62572 15980 62612 17032
rect 62667 17032 62668 17072
rect 62708 17032 62709 17072
rect 62667 17023 62709 17032
rect 62668 16232 62708 17023
rect 62764 16988 62804 17116
rect 62855 17072 62895 17472
rect 63145 17072 63185 17472
rect 63255 17072 63295 17472
rect 63545 17072 63585 17472
rect 63655 17072 63695 17472
rect 63945 17156 63985 17472
rect 62855 17032 63092 17072
rect 63145 17032 63188 17072
rect 62764 16948 62996 16988
rect 62668 16157 62708 16192
rect 62956 16232 62996 16948
rect 63052 16484 63092 17032
rect 63052 16435 63092 16444
rect 63148 16232 63188 17032
rect 63244 17032 63295 17072
rect 63532 17032 63585 17072
rect 63628 17032 63695 17072
rect 63820 17116 63985 17156
rect 63244 16484 63284 17032
rect 63340 16484 63380 16493
rect 63244 16444 63340 16484
rect 63340 16416 63380 16444
rect 63244 16232 63284 16241
rect 63148 16192 63244 16232
rect 62667 16148 62709 16157
rect 62667 16108 62668 16148
rect 62708 16108 62709 16148
rect 62667 16099 62709 16108
rect 62764 16064 62804 16073
rect 62764 15980 62804 16024
rect 62572 15940 62804 15980
rect 62091 15896 62133 15905
rect 62091 15856 62092 15896
rect 62132 15856 62133 15896
rect 62091 15847 62133 15856
rect 61804 15560 61844 15569
rect 61708 15520 61804 15560
rect 61611 15308 61653 15317
rect 61611 15268 61612 15308
rect 61652 15268 61653 15308
rect 61611 15259 61653 15268
rect 60940 14972 60980 14981
rect 60748 14932 60940 14972
rect 60940 14923 60980 14932
rect 61420 14888 61460 14897
rect 61036 14848 61420 14888
rect 60748 14804 60788 14815
rect 61036 14804 61076 14848
rect 61420 14839 61460 14848
rect 60748 14729 60788 14764
rect 60940 14764 61076 14804
rect 61611 14804 61653 14813
rect 61611 14764 61612 14804
rect 61652 14764 61653 14804
rect 60747 14720 60789 14729
rect 60747 14680 60748 14720
rect 60788 14680 60789 14720
rect 60747 14671 60789 14680
rect 60940 14720 60980 14764
rect 61611 14755 61653 14764
rect 60556 14552 60596 14561
rect 60459 14384 60501 14393
rect 60459 14344 60460 14384
rect 60500 14344 60501 14384
rect 60459 14335 60501 14344
rect 60460 12980 60500 14335
rect 60556 13973 60596 14512
rect 60651 14300 60693 14309
rect 60940 14300 60980 14680
rect 60651 14260 60652 14300
rect 60692 14260 60693 14300
rect 60651 14251 60693 14260
rect 60748 14260 60980 14300
rect 61132 14720 61172 14729
rect 60555 13964 60597 13973
rect 60555 13924 60556 13964
rect 60596 13924 60597 13964
rect 60555 13915 60597 13924
rect 60556 13796 60596 13805
rect 60652 13796 60692 14251
rect 60596 13756 60692 13796
rect 60556 13747 60596 13756
rect 60460 12940 60596 12980
rect 60556 11696 60596 12940
rect 60748 11873 60788 14260
rect 61132 14216 61172 14680
rect 61227 14720 61269 14729
rect 61227 14680 61228 14720
rect 61268 14680 61269 14720
rect 61227 14671 61269 14680
rect 61228 14586 61268 14671
rect 61612 14670 61652 14755
rect 61708 14393 61748 15520
rect 61804 15511 61844 15520
rect 61995 15560 62037 15569
rect 62956 15560 62996 16192
rect 61995 15520 61996 15560
rect 62036 15520 62037 15560
rect 61995 15511 62037 15520
rect 62668 15520 62996 15560
rect 61996 14804 62036 15511
rect 62379 15308 62421 15317
rect 62379 15268 62380 15308
rect 62420 15268 62421 15308
rect 62379 15259 62421 15268
rect 61996 14755 62036 14764
rect 62188 14720 62228 14729
rect 62188 14561 62228 14680
rect 62283 14720 62325 14729
rect 62283 14680 62284 14720
rect 62324 14680 62325 14720
rect 62283 14671 62325 14680
rect 62380 14720 62420 15259
rect 62284 14586 62324 14671
rect 61803 14552 61845 14561
rect 61803 14512 61804 14552
rect 61844 14512 61845 14552
rect 61803 14503 61845 14512
rect 62187 14552 62229 14561
rect 62187 14512 62188 14552
rect 62228 14512 62229 14552
rect 62187 14503 62229 14512
rect 61804 14418 61844 14503
rect 61707 14384 61749 14393
rect 61707 14344 61708 14384
rect 61748 14344 61749 14384
rect 61707 14335 61749 14344
rect 60940 14176 61172 14216
rect 60843 14048 60885 14057
rect 60843 14008 60844 14048
rect 60884 14008 60885 14048
rect 60843 13999 60885 14008
rect 60747 11864 60789 11873
rect 60747 11824 60748 11864
rect 60788 11824 60789 11864
rect 60747 11815 60789 11824
rect 60748 11705 60788 11815
rect 60556 11647 60596 11656
rect 60747 11696 60789 11705
rect 60747 11656 60748 11696
rect 60788 11656 60789 11696
rect 60747 11647 60789 11656
rect 60844 11537 60884 13999
rect 60940 13796 60980 14176
rect 62380 14141 62420 14680
rect 62572 14552 62612 14563
rect 62572 14477 62612 14512
rect 62571 14468 62613 14477
rect 62571 14428 62572 14468
rect 62612 14428 62613 14468
rect 62571 14419 62613 14428
rect 62475 14384 62517 14393
rect 62475 14344 62476 14384
rect 62516 14344 62517 14384
rect 62475 14335 62517 14344
rect 61419 14132 61461 14141
rect 61419 14092 61420 14132
rect 61460 14092 61461 14132
rect 61419 14083 61461 14092
rect 62379 14132 62421 14141
rect 62379 14092 62380 14132
rect 62420 14092 62421 14132
rect 62379 14083 62421 14092
rect 60940 12368 60980 13756
rect 61036 14048 61076 14057
rect 61036 13460 61076 14008
rect 61036 13411 61076 13420
rect 61228 14048 61268 14057
rect 61131 13040 61173 13049
rect 61131 13000 61132 13040
rect 61172 13000 61173 13040
rect 61131 12991 61173 13000
rect 61132 12536 61172 12991
rect 61228 12704 61268 14008
rect 61323 13208 61365 13217
rect 61323 13168 61324 13208
rect 61364 13168 61365 13208
rect 61323 13159 61365 13168
rect 61420 13208 61460 14083
rect 62476 14057 62516 14335
rect 61612 14048 61652 14057
rect 61612 13385 61652 14008
rect 62475 14048 62517 14057
rect 62475 14008 62476 14048
rect 62516 14008 62517 14048
rect 62475 13999 62517 14008
rect 61707 13964 61749 13973
rect 61707 13924 61708 13964
rect 61748 13924 61749 13964
rect 61707 13915 61749 13924
rect 61611 13376 61653 13385
rect 61611 13336 61612 13376
rect 61652 13336 61653 13376
rect 61611 13327 61653 13336
rect 61420 13159 61460 13168
rect 61708 13208 61748 13915
rect 62476 13914 62516 13999
rect 62572 13973 62612 14419
rect 62571 13964 62613 13973
rect 62571 13924 62572 13964
rect 62612 13924 62613 13964
rect 62571 13915 62613 13924
rect 62475 13376 62517 13385
rect 62475 13336 62476 13376
rect 62516 13336 62517 13376
rect 62475 13327 62517 13336
rect 61995 13292 62037 13301
rect 61995 13252 61996 13292
rect 62036 13252 62132 13292
rect 61995 13243 62037 13252
rect 61324 13074 61364 13159
rect 61708 12980 61748 13168
rect 62092 13208 62132 13252
rect 62476 13242 62516 13327
rect 62092 13159 62132 13168
rect 62188 13208 62228 13217
rect 61996 13049 62036 13134
rect 61995 13040 62037 13049
rect 61995 13000 61996 13040
rect 62036 13000 62037 13040
rect 61995 12991 62037 13000
rect 61708 12940 61844 12980
rect 62188 12965 62228 13168
rect 62283 13208 62325 13217
rect 62283 13168 62284 13208
rect 62324 13168 62325 13208
rect 62283 13159 62325 13168
rect 62284 13074 62324 13159
rect 61420 12704 61460 12713
rect 61228 12664 61420 12704
rect 61420 12655 61460 12664
rect 61707 12620 61749 12629
rect 61707 12580 61708 12620
rect 61748 12580 61749 12620
rect 61707 12571 61749 12580
rect 61324 12536 61364 12545
rect 61132 12496 61324 12536
rect 61324 12487 61364 12496
rect 61516 12536 61556 12545
rect 61516 12368 61556 12496
rect 61612 12536 61652 12545
rect 61612 12377 61652 12496
rect 60940 12328 61556 12368
rect 61611 12368 61653 12377
rect 61611 12328 61612 12368
rect 61652 12328 61653 12368
rect 61611 12319 61653 12328
rect 61035 11948 61077 11957
rect 61035 11908 61036 11948
rect 61076 11908 61077 11948
rect 61035 11899 61077 11908
rect 61708 11948 61748 12571
rect 61708 11899 61748 11908
rect 60843 11528 60885 11537
rect 60843 11488 60844 11528
rect 60884 11488 60885 11528
rect 60843 11479 60885 11488
rect 60939 11192 60981 11201
rect 60939 11152 60940 11192
rect 60980 11152 60981 11192
rect 60939 11143 60981 11152
rect 60940 11058 60980 11143
rect 60363 10520 60405 10529
rect 60363 10480 60364 10520
rect 60404 10480 60405 10520
rect 60363 10471 60405 10480
rect 60268 10352 60308 10361
rect 60268 10025 60308 10312
rect 60267 10016 60309 10025
rect 60267 9976 60268 10016
rect 60308 9976 60309 10016
rect 60267 9967 60309 9976
rect 60843 9512 60885 9521
rect 60843 9472 60844 9512
rect 60884 9472 60885 9512
rect 60843 9463 60885 9472
rect 60172 9388 60308 9428
rect 59884 9304 60020 9344
rect 59883 9092 59925 9101
rect 59883 9052 59884 9092
rect 59924 9052 59925 9092
rect 59883 9043 59925 9052
rect 59307 8336 59349 8345
rect 59307 8296 59308 8336
rect 59348 8296 59349 8336
rect 59307 8287 59349 8296
rect 59019 8000 59061 8009
rect 59019 7960 59020 8000
rect 59060 7960 59061 8000
rect 59019 7951 59061 7960
rect 58923 7160 58965 7169
rect 58923 7120 58924 7160
rect 58964 7120 58965 7160
rect 58923 7111 58965 7120
rect 58347 6616 58348 6656
rect 58388 6616 58389 6656
rect 58347 6607 58389 6616
rect 58636 6616 58772 6656
rect 58827 6656 58869 6665
rect 58827 6616 58828 6656
rect 58868 6616 58869 6656
rect 58252 6488 58292 6497
rect 58252 6329 58292 6448
rect 58348 6488 58388 6607
rect 58348 6439 58388 6448
rect 58539 6488 58581 6497
rect 58539 6448 58540 6488
rect 58580 6448 58581 6488
rect 58539 6439 58581 6448
rect 58636 6488 58676 6616
rect 58827 6607 58869 6616
rect 58540 6354 58580 6439
rect 58251 6320 58293 6329
rect 58251 6280 58252 6320
rect 58292 6280 58293 6320
rect 58251 6271 58293 6280
rect 58155 5564 58197 5573
rect 58155 5524 58156 5564
rect 58196 5524 58197 5564
rect 58155 5515 58197 5524
rect 57772 4348 57908 4388
rect 57195 4339 57237 4348
rect 56428 4087 56468 4096
rect 56524 4052 56564 4063
rect 56524 3977 56564 4012
rect 56523 3968 56565 3977
rect 56523 3928 56524 3968
rect 56564 3928 56565 3968
rect 56523 3919 56565 3928
rect 56716 3548 56756 4339
rect 56716 3499 56756 3508
rect 56812 4304 56852 4313
rect 56619 3464 56661 3473
rect 56619 3424 56620 3464
rect 56660 3424 56661 3464
rect 56619 3415 56661 3424
rect 56812 3464 56852 4264
rect 57003 4136 57045 4145
rect 57003 4096 57004 4136
rect 57044 4096 57045 4136
rect 57003 4087 57045 4096
rect 57196 4136 57236 4339
rect 57291 4304 57333 4313
rect 57291 4264 57292 4304
rect 57332 4264 57333 4304
rect 57291 4255 57333 4264
rect 57196 4087 57236 4096
rect 57292 4136 57332 4255
rect 57868 4136 57908 4348
rect 57964 4313 58004 4398
rect 57963 4304 58005 4313
rect 57963 4264 57964 4304
rect 58004 4264 58005 4304
rect 57963 4255 58005 4264
rect 57964 4136 58004 4145
rect 57868 4096 57964 4136
rect 57292 4087 57332 4096
rect 57964 4087 58004 4096
rect 58156 4136 58196 5515
rect 58539 4724 58581 4733
rect 58539 4684 58540 4724
rect 58580 4684 58581 4724
rect 58539 4675 58581 4684
rect 58540 4590 58580 4675
rect 58636 4229 58676 6448
rect 58732 6488 58772 6499
rect 58732 6413 58772 6448
rect 58827 6488 58869 6497
rect 58827 6448 58828 6488
rect 58868 6448 58869 6488
rect 58827 6439 58869 6448
rect 58731 6404 58773 6413
rect 58731 6364 58732 6404
rect 58772 6364 58773 6404
rect 58731 6355 58773 6364
rect 58828 6354 58868 6439
rect 58827 5480 58869 5489
rect 58827 5440 58828 5480
rect 58868 5440 58869 5480
rect 58827 5431 58869 5440
rect 58828 5060 58868 5431
rect 58828 5011 58868 5020
rect 58924 4892 58964 7111
rect 59020 6833 59060 7951
rect 59211 7076 59253 7085
rect 59211 7036 59212 7076
rect 59252 7036 59253 7076
rect 59211 7027 59253 7036
rect 59212 6992 59252 7027
rect 59019 6824 59061 6833
rect 59019 6784 59020 6824
rect 59060 6784 59061 6824
rect 59019 6775 59061 6784
rect 59019 6656 59061 6665
rect 59019 6616 59020 6656
rect 59060 6616 59061 6656
rect 59019 6607 59061 6616
rect 59020 6413 59060 6607
rect 59212 6497 59252 6952
rect 59308 6656 59348 8287
rect 59691 7244 59733 7253
rect 59691 7204 59692 7244
rect 59732 7204 59733 7244
rect 59691 7195 59733 7204
rect 59692 7160 59732 7195
rect 59692 7109 59732 7120
rect 59691 6740 59733 6749
rect 59691 6700 59692 6740
rect 59732 6700 59733 6740
rect 59691 6691 59733 6700
rect 59308 6616 59636 6656
rect 59211 6488 59253 6497
rect 59211 6448 59212 6488
rect 59252 6448 59253 6488
rect 59211 6439 59253 6448
rect 59308 6488 59348 6616
rect 59308 6439 59348 6448
rect 59499 6488 59541 6497
rect 59499 6448 59500 6488
rect 59540 6448 59541 6488
rect 59499 6439 59541 6448
rect 59019 6404 59061 6413
rect 59019 6364 59020 6404
rect 59060 6364 59061 6404
rect 59019 6355 59061 6364
rect 58828 4852 58964 4892
rect 58635 4220 58677 4229
rect 58635 4180 58636 4220
rect 58676 4180 58677 4220
rect 58635 4171 58677 4180
rect 58156 4087 58196 4096
rect 58251 4136 58293 4145
rect 58251 4096 58252 4136
rect 58292 4096 58293 4136
rect 58251 4087 58293 4096
rect 57004 4002 57044 4087
rect 58252 4002 58292 4087
rect 57100 3968 57140 3977
rect 57100 3557 57140 3928
rect 58828 3884 58868 4852
rect 58923 4136 58965 4145
rect 58923 4096 58924 4136
rect 58964 4096 58965 4136
rect 58923 4087 58965 4096
rect 59020 4136 59060 6355
rect 59212 6354 59252 6439
rect 59500 6354 59540 6439
rect 59500 6236 59540 6245
rect 59212 5648 59252 5657
rect 59212 5144 59252 5608
rect 59403 5648 59445 5657
rect 59403 5608 59404 5648
rect 59444 5608 59445 5648
rect 59403 5599 59445 5608
rect 59500 5648 59540 6196
rect 59500 5599 59540 5608
rect 59404 5514 59444 5599
rect 59307 5480 59349 5489
rect 59307 5440 59308 5480
rect 59348 5440 59349 5480
rect 59307 5431 59349 5440
rect 59308 5346 59348 5431
rect 59212 5104 59348 5144
rect 59211 4976 59253 4985
rect 59211 4936 59212 4976
rect 59252 4936 59253 4976
rect 59211 4927 59253 4936
rect 59212 4842 59252 4927
rect 59115 4220 59157 4229
rect 59115 4180 59116 4220
rect 59156 4180 59157 4220
rect 59115 4171 59157 4180
rect 58924 4002 58964 4087
rect 58828 3844 58964 3884
rect 57099 3548 57141 3557
rect 57099 3508 57100 3548
rect 57140 3508 57141 3548
rect 57099 3499 57141 3508
rect 56812 3415 56852 3424
rect 58827 3464 58869 3473
rect 58827 3424 58828 3464
rect 58868 3424 58869 3464
rect 58827 3415 58869 3424
rect 56620 2900 56660 3415
rect 56620 2860 56852 2900
rect 56523 2792 56565 2801
rect 56523 2752 56524 2792
rect 56564 2752 56565 2792
rect 56523 2743 56565 2752
rect 56332 2575 56372 2584
rect 56524 2624 56564 2743
rect 56524 2575 56564 2584
rect 56620 2624 56660 2633
rect 56812 2624 56852 2860
rect 58828 2876 58868 3415
rect 58924 2885 58964 3844
rect 59020 3137 59060 4096
rect 59116 4136 59156 4171
rect 59116 4085 59156 4096
rect 59212 4136 59252 4145
rect 59308 4136 59348 5104
rect 59596 4313 59636 6616
rect 59692 6581 59732 6691
rect 59691 6572 59733 6581
rect 59691 6532 59692 6572
rect 59732 6532 59733 6572
rect 59691 6523 59733 6532
rect 59788 6497 59828 8632
rect 59787 6488 59829 6497
rect 59787 6448 59788 6488
rect 59828 6448 59829 6488
rect 59787 6439 59829 6448
rect 59692 5816 59732 5825
rect 59692 4985 59732 5776
rect 59691 4976 59733 4985
rect 59691 4936 59692 4976
rect 59732 4936 59733 4976
rect 59691 4927 59733 4936
rect 59403 4304 59445 4313
rect 59403 4264 59404 4304
rect 59444 4264 59445 4304
rect 59403 4255 59445 4264
rect 59595 4304 59637 4313
rect 59595 4264 59596 4304
rect 59636 4264 59637 4304
rect 59595 4255 59637 4264
rect 59252 4096 59348 4136
rect 59212 4087 59252 4096
rect 59308 3464 59348 3473
rect 59404 3464 59444 4255
rect 59499 3716 59541 3725
rect 59499 3676 59500 3716
rect 59540 3676 59541 3716
rect 59499 3667 59541 3676
rect 59348 3424 59444 3464
rect 59500 3464 59540 3667
rect 59308 3415 59348 3424
rect 59404 3212 59444 3221
rect 59116 3172 59404 3212
rect 59019 3128 59061 3137
rect 59019 3088 59020 3128
rect 59060 3088 59061 3128
rect 59019 3079 59061 3088
rect 58828 2827 58868 2836
rect 58923 2876 58965 2885
rect 58923 2836 58924 2876
rect 58964 2836 58965 2876
rect 58923 2827 58965 2836
rect 56907 2792 56949 2801
rect 56907 2752 56908 2792
rect 56948 2752 56949 2792
rect 56907 2743 56949 2752
rect 56908 2658 56948 2743
rect 57291 2708 57333 2717
rect 57291 2668 57292 2708
rect 57332 2668 57333 2708
rect 57291 2659 57333 2668
rect 58731 2708 58773 2717
rect 58731 2668 58732 2708
rect 58772 2668 58773 2708
rect 58731 2659 58773 2668
rect 56660 2584 56756 2624
rect 56620 2575 56660 2584
rect 56428 2456 56468 2465
rect 56468 2416 56660 2456
rect 56428 2407 56468 2416
rect 56523 2120 56565 2129
rect 56523 2080 56524 2120
rect 56564 2080 56565 2120
rect 56523 2071 56565 2080
rect 56236 1903 56276 1912
rect 56331 1952 56373 1961
rect 56331 1912 56332 1952
rect 56372 1912 56373 1952
rect 56331 1903 56373 1912
rect 56332 1818 56372 1903
rect 56524 1205 56564 2071
rect 56620 2036 56660 2416
rect 56620 1987 56660 1996
rect 56523 1196 56565 1205
rect 56523 1156 56524 1196
rect 56564 1156 56565 1196
rect 56716 1196 56756 2584
rect 56812 2575 56852 2584
rect 57004 2624 57044 2633
rect 57004 2372 57044 2584
rect 56812 2332 57044 2372
rect 57196 2624 57236 2633
rect 56812 1364 56852 2332
rect 57196 2129 57236 2584
rect 57292 2624 57332 2659
rect 57195 2120 57237 2129
rect 57195 2080 57196 2120
rect 57236 2080 57237 2120
rect 57195 2071 57237 2080
rect 57003 1952 57045 1961
rect 57003 1912 57004 1952
rect 57044 1912 57045 1952
rect 57003 1903 57045 1912
rect 57004 1818 57044 1903
rect 57195 1448 57237 1457
rect 57195 1408 57196 1448
rect 57236 1408 57237 1448
rect 57195 1399 57237 1408
rect 56812 1315 56852 1324
rect 57100 1280 57140 1289
rect 56908 1240 57100 1280
rect 56908 1196 56948 1240
rect 57100 1231 57140 1240
rect 56716 1156 56948 1196
rect 56523 1147 56565 1156
rect 56140 1063 56180 1072
rect 56427 1112 56469 1121
rect 56427 1072 56428 1112
rect 56468 1072 56469 1112
rect 56427 1063 56469 1072
rect 56524 1112 56564 1147
rect 57196 1121 57236 1399
rect 56428 978 56468 1063
rect 56524 1062 56564 1072
rect 57004 1112 57044 1121
rect 57004 860 57044 1072
rect 57195 1112 57237 1121
rect 57195 1072 57196 1112
rect 57236 1072 57237 1112
rect 57195 1063 57237 1072
rect 57196 978 57236 1063
rect 57292 860 57332 2584
rect 57484 2624 57524 2633
rect 57484 2540 57524 2584
rect 57579 2540 57621 2549
rect 57484 2500 57580 2540
rect 57620 2500 57621 2540
rect 57579 2491 57621 2500
rect 57388 2456 57428 2465
rect 57428 2416 57524 2456
rect 57388 2407 57428 2416
rect 57387 1952 57429 1961
rect 57387 1912 57388 1952
rect 57428 1912 57429 1952
rect 57387 1903 57429 1912
rect 57388 1280 57428 1903
rect 57388 1231 57428 1240
rect 57484 1121 57524 2416
rect 57867 1952 57909 1961
rect 57867 1912 57868 1952
rect 57908 1912 57909 1952
rect 57867 1903 57909 1912
rect 57868 1818 57908 1903
rect 57483 1112 57525 1121
rect 57483 1072 57484 1112
rect 57524 1072 57525 1112
rect 57483 1063 57525 1072
rect 58635 1112 58677 1121
rect 58635 1072 58636 1112
rect 58676 1072 58677 1112
rect 58635 1063 58677 1072
rect 58732 1112 58772 2659
rect 58828 2624 58868 2633
rect 58924 2624 58964 2827
rect 59019 2708 59061 2717
rect 59019 2668 59020 2708
rect 59060 2668 59061 2708
rect 59019 2659 59061 2668
rect 58868 2584 58964 2624
rect 59020 2624 59060 2659
rect 58828 2575 58868 2584
rect 59020 2573 59060 2584
rect 59116 2624 59156 3172
rect 59404 3163 59444 3172
rect 59403 3044 59445 3053
rect 59403 3004 59404 3044
rect 59444 3004 59445 3044
rect 59403 2995 59445 3004
rect 59116 2575 59156 2584
rect 59404 2624 59444 2995
rect 59500 2624 59540 3424
rect 59691 3464 59733 3473
rect 59691 3424 59692 3464
rect 59732 3424 59733 3464
rect 59691 3415 59733 3424
rect 59692 3330 59732 3415
rect 59692 2624 59732 2633
rect 59500 2584 59692 2624
rect 59404 2575 59444 2584
rect 59692 2575 59732 2584
rect 59787 2540 59829 2549
rect 59787 2500 59788 2540
rect 59828 2500 59829 2540
rect 59787 2491 59829 2500
rect 59788 2406 59828 2491
rect 59115 1952 59157 1961
rect 59115 1912 59116 1952
rect 59156 1912 59157 1952
rect 59115 1903 59157 1912
rect 59212 1952 59252 1961
rect 59019 1700 59061 1709
rect 59019 1660 59020 1700
rect 59060 1660 59061 1700
rect 59019 1651 59061 1660
rect 59020 1457 59060 1651
rect 59019 1448 59061 1457
rect 59019 1408 59020 1448
rect 59060 1408 59061 1448
rect 59019 1399 59061 1408
rect 58923 1364 58965 1373
rect 58923 1324 58924 1364
rect 58964 1324 58965 1364
rect 58923 1315 58965 1324
rect 58924 1230 58964 1315
rect 58732 1063 58772 1072
rect 58924 1112 58964 1121
rect 58636 978 58676 1063
rect 58924 953 58964 1072
rect 59116 1112 59156 1903
rect 59212 1373 59252 1912
rect 59596 1952 59636 1961
rect 59211 1364 59253 1373
rect 59211 1324 59212 1364
rect 59252 1324 59253 1364
rect 59211 1315 59253 1324
rect 59596 1289 59636 1912
rect 59595 1280 59637 1289
rect 59595 1240 59596 1280
rect 59636 1240 59637 1280
rect 59595 1231 59637 1240
rect 59884 1121 59924 9043
rect 59980 8672 60020 9304
rect 60171 9260 60213 9269
rect 60171 9220 60172 9260
rect 60212 9220 60213 9260
rect 60171 9211 60213 9220
rect 59980 8345 60020 8632
rect 60075 8672 60117 8681
rect 60075 8632 60076 8672
rect 60116 8632 60117 8672
rect 60075 8623 60117 8632
rect 60172 8672 60212 9211
rect 60172 8623 60212 8632
rect 60076 8538 60116 8623
rect 60268 8513 60308 9388
rect 60844 9378 60884 9463
rect 60363 9176 60405 9185
rect 60363 9136 60364 9176
rect 60404 9136 60405 9176
rect 60363 9127 60405 9136
rect 60267 8504 60309 8513
rect 60267 8464 60268 8504
rect 60308 8464 60309 8504
rect 60267 8455 60309 8464
rect 59979 8336 60021 8345
rect 59979 8296 59980 8336
rect 60020 8296 60308 8336
rect 59979 8287 60021 8296
rect 59980 8202 60020 8287
rect 60075 8168 60117 8177
rect 60075 8128 60076 8168
rect 60116 8128 60117 8168
rect 60075 8119 60117 8128
rect 60076 8000 60116 8119
rect 59980 7960 60076 8000
rect 59980 7160 60020 7960
rect 60076 7951 60116 7960
rect 60268 8000 60308 8296
rect 60268 7951 60308 7960
rect 60364 7841 60404 9127
rect 60940 8840 60980 8849
rect 60460 8000 60500 8009
rect 60844 8000 60884 8009
rect 60940 8000 60980 8800
rect 60500 7960 60788 8000
rect 60460 7951 60500 7960
rect 60363 7832 60405 7841
rect 60363 7792 60364 7832
rect 60404 7792 60405 7832
rect 60363 7783 60405 7792
rect 60171 7748 60213 7757
rect 60171 7708 60172 7748
rect 60212 7708 60213 7748
rect 60171 7699 60213 7708
rect 60172 7614 60212 7699
rect 60364 7244 60404 7783
rect 60555 7748 60597 7757
rect 60555 7708 60556 7748
rect 60596 7708 60597 7748
rect 60555 7699 60597 7708
rect 60459 7244 60501 7253
rect 60364 7204 60460 7244
rect 60500 7204 60501 7244
rect 60459 7195 60501 7204
rect 59980 7111 60020 7120
rect 60075 7076 60117 7085
rect 60075 7036 60076 7076
rect 60116 7036 60117 7076
rect 60075 7027 60117 7036
rect 60076 6942 60116 7027
rect 60364 6950 60404 6959
rect 60171 6488 60213 6497
rect 60171 6448 60172 6488
rect 60212 6448 60213 6488
rect 60171 6439 60213 6448
rect 60364 6488 60404 6910
rect 60364 6439 60404 6448
rect 60075 5732 60117 5741
rect 60075 5692 60076 5732
rect 60116 5692 60117 5732
rect 60075 5683 60117 5692
rect 60076 4985 60116 5683
rect 60172 5069 60212 6439
rect 60267 6320 60309 6329
rect 60267 6280 60268 6320
rect 60308 6280 60309 6320
rect 60267 6271 60309 6280
rect 60268 6186 60308 6271
rect 60364 5648 60404 5657
rect 60460 5648 60500 7195
rect 60556 7160 60596 7699
rect 60556 7111 60596 7120
rect 60652 7160 60692 7169
rect 60652 6329 60692 7120
rect 60748 7076 60788 7960
rect 60884 7960 60980 8000
rect 60844 7951 60884 7960
rect 61036 7328 61076 11899
rect 61804 11453 61844 12940
rect 62187 12956 62229 12965
rect 62187 12916 62188 12956
rect 62228 12916 62229 12956
rect 62187 12907 62229 12916
rect 62091 12704 62133 12713
rect 62091 12664 62092 12704
rect 62132 12664 62133 12704
rect 62091 12655 62133 12664
rect 62092 12536 62132 12655
rect 61996 12496 62092 12536
rect 61803 11444 61845 11453
rect 61803 11404 61804 11444
rect 61844 11404 61845 11444
rect 61803 11395 61845 11404
rect 61804 11033 61844 11395
rect 61803 11024 61845 11033
rect 61803 10984 61804 11024
rect 61844 10984 61845 11024
rect 61803 10975 61845 10984
rect 61996 10361 62036 12496
rect 62092 12487 62132 12496
rect 62284 12536 62324 12547
rect 62284 12461 62324 12496
rect 62380 12536 62420 12545
rect 62283 12452 62325 12461
rect 62283 12412 62284 12452
rect 62324 12412 62325 12452
rect 62283 12403 62325 12412
rect 62091 12368 62133 12377
rect 62091 12328 62092 12368
rect 62132 12328 62133 12368
rect 62091 12319 62133 12328
rect 62092 12234 62132 12319
rect 62092 11864 62132 11873
rect 62132 11824 62228 11864
rect 62092 11815 62132 11824
rect 62091 11696 62133 11705
rect 62091 11656 62092 11696
rect 62132 11656 62133 11696
rect 62091 11647 62133 11656
rect 62092 11024 62132 11647
rect 62188 11033 62228 11824
rect 62380 11201 62420 12496
rect 62571 11948 62613 11957
rect 62571 11908 62572 11948
rect 62612 11908 62613 11948
rect 62571 11899 62613 11908
rect 62572 11789 62612 11899
rect 62571 11780 62613 11789
rect 62571 11740 62572 11780
rect 62612 11740 62613 11780
rect 62571 11731 62613 11740
rect 62379 11192 62421 11201
rect 62379 11152 62380 11192
rect 62420 11152 62421 11192
rect 62379 11143 62421 11152
rect 62092 10975 62132 10984
rect 62187 11024 62229 11033
rect 62187 10984 62188 11024
rect 62228 10984 62229 11024
rect 62187 10975 62229 10984
rect 61995 10352 62037 10361
rect 61995 10312 61996 10352
rect 62036 10312 62037 10352
rect 61995 10303 62037 10312
rect 62380 10352 62420 10361
rect 61995 9680 62037 9689
rect 61995 9640 61996 9680
rect 62036 9640 62037 9680
rect 61995 9631 62037 9640
rect 61996 9546 62036 9631
rect 62187 9596 62229 9605
rect 62187 9556 62188 9596
rect 62228 9556 62229 9596
rect 62187 9547 62229 9556
rect 62188 9462 62228 9547
rect 62380 9512 62420 10312
rect 62572 9512 62612 9521
rect 62380 9472 62572 9512
rect 62572 9463 62612 9472
rect 61995 9260 62037 9269
rect 61995 9220 61996 9260
rect 62036 9220 62037 9260
rect 61995 9211 62037 9220
rect 61996 9126 62036 9211
rect 62668 9017 62708 15520
rect 63244 15476 63284 16192
rect 63532 16232 63572 17032
rect 63628 16484 63668 17032
rect 63628 16435 63668 16444
rect 63532 16073 63572 16192
rect 63820 16232 63860 17116
rect 64055 17072 64095 17472
rect 64345 17156 64385 17472
rect 63916 17032 64095 17072
rect 64300 17116 64385 17156
rect 63916 16484 63956 17032
rect 63916 16435 63956 16444
rect 63531 16064 63573 16073
rect 63531 16024 63532 16064
rect 63572 16024 63573 16064
rect 63531 16015 63573 16024
rect 63820 15728 63860 16192
rect 62860 15436 63284 15476
rect 63532 15688 63860 15728
rect 64108 16232 64148 16241
rect 64300 16232 64340 17116
rect 64455 17072 64495 17472
rect 64587 17156 64629 17165
rect 64745 17156 64785 17472
rect 64855 17165 64895 17472
rect 64587 17116 64588 17156
rect 64628 17116 64629 17156
rect 64587 17107 64629 17116
rect 64684 17116 64785 17156
rect 64854 17156 64896 17165
rect 65145 17156 65185 17472
rect 64854 17116 64855 17156
rect 64895 17116 64896 17156
rect 64148 16192 64340 16232
rect 64396 17032 64495 17072
rect 62763 14888 62805 14897
rect 62763 14848 62764 14888
rect 62804 14848 62805 14888
rect 62763 14839 62805 14848
rect 62764 14804 62804 14839
rect 62764 14753 62804 14764
rect 62860 14636 62900 15436
rect 62955 15308 62997 15317
rect 62955 15268 62956 15308
rect 62996 15268 62997 15308
rect 62955 15259 62997 15268
rect 62956 15174 62996 15259
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 62764 14596 62900 14636
rect 62764 12209 62804 14596
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 63532 13469 63572 15688
rect 64108 15401 64148 16192
rect 64204 16064 64244 16073
rect 64396 16064 64436 17032
rect 64588 16484 64628 17107
rect 64684 16913 64724 17116
rect 64854 17107 64896 17116
rect 64972 17116 65185 17156
rect 64683 16904 64725 16913
rect 64683 16864 64684 16904
rect 64724 16864 64725 16904
rect 64683 16855 64725 16864
rect 64588 16435 64628 16444
rect 64492 16232 64532 16241
rect 64684 16232 64724 16855
rect 64972 16241 65012 17116
rect 65255 17072 65295 17472
rect 65545 17156 65585 17472
rect 65068 17032 65295 17072
rect 65356 17116 65585 17156
rect 65068 16484 65108 17032
rect 65356 16577 65396 17116
rect 65655 17072 65695 17472
rect 65945 17156 65985 17472
rect 65452 17032 65695 17072
rect 65740 17116 65985 17156
rect 65355 16568 65397 16577
rect 65355 16528 65356 16568
rect 65396 16528 65397 16568
rect 65355 16519 65397 16528
rect 65068 16435 65108 16444
rect 64532 16192 64724 16232
rect 64971 16232 65013 16241
rect 64971 16192 64972 16232
rect 65012 16192 65013 16232
rect 64492 16183 64532 16192
rect 64971 16183 65013 16192
rect 65356 16232 65396 16519
rect 65452 16484 65492 17032
rect 65452 16435 65492 16444
rect 65356 16183 65396 16192
rect 65740 16232 65780 17116
rect 66055 17072 66095 17472
rect 66345 17156 66385 17472
rect 65836 17032 66095 17072
rect 66316 17116 66385 17156
rect 65836 16484 65876 17032
rect 65836 16435 65876 16444
rect 64972 16098 65012 16183
rect 64244 16024 64436 16064
rect 64204 16015 64244 16024
rect 64491 15728 64533 15737
rect 64491 15688 64492 15728
rect 64532 15688 64533 15728
rect 64491 15679 64533 15688
rect 64779 15728 64821 15737
rect 64779 15688 64780 15728
rect 64820 15688 64821 15728
rect 64779 15679 64821 15688
rect 64107 15392 64149 15401
rect 64107 15352 64108 15392
rect 64148 15352 64149 15392
rect 64107 15343 64149 15352
rect 64108 14888 64148 14897
rect 63916 14848 64108 14888
rect 63724 14720 63764 14729
rect 63724 14393 63764 14680
rect 63819 14720 63861 14729
rect 63819 14680 63820 14720
rect 63860 14680 63861 14720
rect 63819 14671 63861 14680
rect 63916 14720 63956 14848
rect 64108 14839 64148 14848
rect 63916 14671 63956 14680
rect 64492 14720 64532 15679
rect 64780 15560 64820 15679
rect 64780 15511 64820 15520
rect 64971 15560 65013 15569
rect 64971 15520 64972 15560
rect 65012 15520 65013 15560
rect 64971 15511 65013 15520
rect 65452 15560 65492 15569
rect 64972 15426 65012 15511
rect 64876 15308 64916 15317
rect 64916 15268 65108 15308
rect 64876 15259 64916 15268
rect 64492 14671 64532 14680
rect 64683 14720 64725 14729
rect 64683 14680 64684 14720
rect 64724 14680 64725 14720
rect 64683 14671 64725 14680
rect 64780 14720 64820 14729
rect 65068 14720 65108 15268
rect 65356 14972 65396 14981
rect 65452 14972 65492 15520
rect 65740 15317 65780 16192
rect 66124 16232 66164 16241
rect 66316 16232 66356 17116
rect 66455 17072 66495 17472
rect 66603 17156 66645 17165
rect 66745 17156 66785 17472
rect 66855 17165 66895 17472
rect 66603 17116 66604 17156
rect 66644 17116 66645 17156
rect 66603 17107 66645 17116
rect 66700 17116 66785 17156
rect 66854 17156 66896 17165
rect 67145 17156 67185 17472
rect 66854 17116 66855 17156
rect 66895 17116 66896 17156
rect 66164 16192 66356 16232
rect 66412 17032 66495 17072
rect 66124 15989 66164 16192
rect 66220 16064 66260 16073
rect 66412 16064 66452 17032
rect 66604 16484 66644 17107
rect 66604 16435 66644 16444
rect 66260 16024 66452 16064
rect 66508 16232 66548 16241
rect 66700 16232 66740 17116
rect 66854 17107 66896 17116
rect 66988 17116 67185 17156
rect 66548 16192 66740 16232
rect 66795 16232 66837 16241
rect 66988 16232 67028 17116
rect 67255 17072 67295 17472
rect 67545 17072 67585 17472
rect 67084 17032 67295 17072
rect 67372 17032 67585 17072
rect 67655 17072 67695 17472
rect 67945 17156 67985 17472
rect 67756 17116 67985 17156
rect 67655 17032 67700 17072
rect 67084 16484 67124 17032
rect 67084 16435 67124 16444
rect 67372 16241 67412 17032
rect 67468 16484 67508 16493
rect 67660 16484 67700 17032
rect 67508 16444 67700 16484
rect 67468 16435 67508 16444
rect 66795 16192 66796 16232
rect 66836 16192 66837 16232
rect 66220 16015 66260 16024
rect 66123 15980 66165 15989
rect 66123 15940 66124 15980
rect 66164 15940 66165 15980
rect 66123 15931 66165 15940
rect 65836 15560 65876 15569
rect 65739 15308 65781 15317
rect 65739 15268 65740 15308
rect 65780 15268 65781 15308
rect 65739 15259 65781 15268
rect 65396 14932 65492 14972
rect 65356 14923 65396 14932
rect 65836 14888 65876 15520
rect 66219 15476 66261 15485
rect 66219 15436 66220 15476
rect 66260 15436 66261 15476
rect 66219 15427 66261 15436
rect 65932 14888 65972 14897
rect 65836 14848 65932 14888
rect 65932 14839 65972 14848
rect 64820 14680 64916 14720
rect 64780 14671 64820 14680
rect 63820 14586 63860 14671
rect 64396 14636 64436 14645
rect 64204 14596 64396 14636
rect 63915 14552 63957 14561
rect 63915 14512 63916 14552
rect 63956 14512 63957 14552
rect 63915 14503 63957 14512
rect 63723 14384 63765 14393
rect 63723 14344 63724 14384
rect 63764 14344 63765 14384
rect 63723 14335 63765 14344
rect 63820 14048 63860 14057
rect 63628 13796 63668 13805
rect 63820 13796 63860 14008
rect 63916 14048 63956 14503
rect 64204 14216 64244 14596
rect 64396 14587 64436 14596
rect 64684 14552 64724 14671
rect 64684 14512 64820 14552
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 64780 14216 64820 14512
rect 64204 14176 64436 14216
rect 64108 14048 64148 14057
rect 63916 13973 63956 14008
rect 64012 14008 64108 14048
rect 63915 13964 63957 13973
rect 63915 13924 63916 13964
rect 63956 13924 63957 13964
rect 63915 13915 63957 13924
rect 63668 13756 63860 13796
rect 63531 13460 63573 13469
rect 63531 13420 63532 13460
rect 63572 13420 63573 13460
rect 63531 13411 63573 13420
rect 62859 13292 62901 13301
rect 62859 13252 62860 13292
rect 62900 13252 62901 13292
rect 62859 13243 62901 13252
rect 62860 13133 62900 13243
rect 63628 13217 63668 13756
rect 64012 13544 64052 14008
rect 64108 13999 64148 14008
rect 64396 13973 64436 14176
rect 64492 14176 64820 14216
rect 64395 13964 64437 13973
rect 64395 13924 64396 13964
rect 64436 13924 64437 13964
rect 64395 13915 64437 13924
rect 64108 13796 64148 13805
rect 64148 13756 64340 13796
rect 64108 13747 64148 13756
rect 64012 13504 64244 13544
rect 64107 13376 64149 13385
rect 64107 13336 64108 13376
rect 64148 13336 64149 13376
rect 64107 13327 64149 13336
rect 63627 13208 63669 13217
rect 63627 13168 63628 13208
rect 63668 13168 63669 13208
rect 63627 13159 63669 13168
rect 63915 13208 63957 13217
rect 63915 13168 63916 13208
rect 63956 13168 63957 13208
rect 63915 13159 63957 13168
rect 64012 13208 64052 13217
rect 62859 13124 62901 13133
rect 62859 13084 62860 13124
rect 62900 13084 62901 13124
rect 62859 13075 62901 13084
rect 62763 12200 62805 12209
rect 62763 12160 62764 12200
rect 62804 12160 62805 12200
rect 62763 12151 62805 12160
rect 62763 11948 62805 11957
rect 62763 11908 62764 11948
rect 62804 11908 62805 11948
rect 62763 11899 62805 11908
rect 62764 11780 62804 11899
rect 62860 11864 62900 13075
rect 63820 13049 63860 13134
rect 63916 13074 63956 13159
rect 63819 13040 63861 13049
rect 63819 13000 63820 13040
rect 63860 13000 63861 13040
rect 63819 12991 63861 13000
rect 64012 12965 64052 13168
rect 64108 13208 64148 13327
rect 64108 13159 64148 13168
rect 63531 12956 63573 12965
rect 63531 12916 63532 12956
rect 63572 12916 63573 12956
rect 63531 12907 63573 12916
rect 64011 12956 64053 12965
rect 64011 12916 64012 12956
rect 64052 12916 64053 12956
rect 64011 12907 64053 12916
rect 63052 12536 63092 12545
rect 62956 12496 63052 12536
rect 62956 11948 62996 12496
rect 63052 12487 63092 12496
rect 63244 12536 63284 12545
rect 63052 12293 63092 12378
rect 63244 12377 63284 12496
rect 63339 12536 63381 12545
rect 63339 12496 63340 12536
rect 63380 12496 63381 12536
rect 63339 12487 63381 12496
rect 63340 12402 63380 12487
rect 63243 12368 63285 12377
rect 63243 12328 63244 12368
rect 63284 12328 63285 12368
rect 63243 12319 63285 12328
rect 63051 12284 63093 12293
rect 63051 12244 63052 12284
rect 63092 12244 63093 12284
rect 63051 12235 63093 12244
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 63532 11957 63572 12907
rect 64204 12713 64244 13504
rect 64300 13208 64340 13756
rect 64396 13385 64436 13915
rect 64395 13376 64437 13385
rect 64395 13336 64396 13376
rect 64436 13336 64437 13376
rect 64395 13327 64437 13336
rect 64300 13159 64340 13168
rect 64396 13208 64436 13217
rect 64492 13208 64532 14176
rect 64684 14048 64724 14057
rect 64588 13460 64628 13469
rect 64684 13460 64724 14008
rect 64628 13420 64724 13460
rect 64588 13411 64628 13420
rect 64436 13168 64532 13208
rect 64588 13208 64628 13217
rect 64396 13159 64436 13168
rect 64588 13049 64628 13168
rect 64587 13040 64629 13049
rect 64587 13000 64588 13040
rect 64628 13000 64629 13040
rect 64587 12991 64629 13000
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 64203 12704 64245 12713
rect 64203 12664 64204 12704
rect 64244 12664 64245 12704
rect 64203 12655 64245 12664
rect 64395 12536 64437 12545
rect 64395 12496 64396 12536
rect 64436 12496 64437 12536
rect 64395 12487 64437 12496
rect 64588 12536 64628 12547
rect 63723 12452 63765 12461
rect 63723 12412 63724 12452
rect 63764 12412 63765 12452
rect 63723 12403 63765 12412
rect 63627 12284 63669 12293
rect 63627 12244 63628 12284
rect 63668 12244 63669 12284
rect 63627 12235 63669 12244
rect 63243 11948 63285 11957
rect 62956 11908 63092 11948
rect 62860 11824 62996 11864
rect 62764 11740 62900 11780
rect 62860 11696 62900 11740
rect 62764 11675 62804 11684
rect 62860 11647 62900 11656
rect 62956 11696 62996 11824
rect 62764 11621 62804 11635
rect 62763 11612 62805 11621
rect 62763 11572 62764 11612
rect 62804 11572 62805 11612
rect 62763 11563 62805 11572
rect 62764 11201 62804 11563
rect 62956 11276 62996 11656
rect 63052 11696 63092 11908
rect 63243 11908 63244 11948
rect 63284 11908 63285 11948
rect 63243 11899 63285 11908
rect 63531 11948 63573 11957
rect 63531 11908 63532 11948
rect 63572 11908 63573 11948
rect 63531 11899 63573 11908
rect 63052 11647 63092 11656
rect 63244 11369 63284 11899
rect 63435 11864 63477 11873
rect 63435 11824 63436 11864
rect 63476 11824 63477 11864
rect 63435 11815 63477 11824
rect 63436 11696 63476 11815
rect 63436 11453 63476 11656
rect 63435 11444 63477 11453
rect 63435 11404 63436 11444
rect 63476 11404 63477 11444
rect 63435 11395 63477 11404
rect 63243 11360 63285 11369
rect 63243 11320 63244 11360
rect 63284 11320 63285 11360
rect 63243 11311 63285 11320
rect 62860 11236 62996 11276
rect 62763 11192 62805 11201
rect 62763 11152 62764 11192
rect 62804 11152 62805 11192
rect 62763 11143 62805 11152
rect 62667 9008 62709 9017
rect 62667 8968 62668 9008
rect 62708 8968 62709 9008
rect 62667 8959 62709 8968
rect 62860 8849 62900 11236
rect 62956 11033 62996 11118
rect 63340 11108 63380 11117
rect 63628 11108 63668 12235
rect 63724 11864 63764 12403
rect 64396 12402 64436 12487
rect 64588 12461 64628 12496
rect 64780 12536 64820 12545
rect 64587 12452 64629 12461
rect 64587 12412 64588 12452
rect 64628 12412 64629 12452
rect 64587 12403 64629 12412
rect 64011 12368 64053 12377
rect 64011 12328 64012 12368
rect 64052 12328 64053 12368
rect 64011 12319 64053 12328
rect 63721 11824 63764 11864
rect 63721 11738 63761 11824
rect 63721 11698 63764 11738
rect 63724 11696 63764 11698
rect 63724 11647 63764 11656
rect 63819 11612 63861 11621
rect 63819 11572 63820 11612
rect 63860 11572 63861 11612
rect 63819 11563 63861 11572
rect 63820 11478 63860 11563
rect 63915 11444 63957 11453
rect 63915 11404 63916 11444
rect 63956 11404 63957 11444
rect 63915 11395 63957 11404
rect 63819 11360 63861 11369
rect 63819 11320 63820 11360
rect 63860 11320 63861 11360
rect 63819 11311 63861 11320
rect 63380 11068 63668 11108
rect 63340 11059 63380 11068
rect 62955 11024 62997 11033
rect 62955 10984 62956 11024
rect 62996 10984 62997 11024
rect 62955 10975 62997 10984
rect 63820 10772 63860 11311
rect 63916 11033 63956 11395
rect 64012 11108 64052 12319
rect 64492 12284 64532 12293
rect 64300 12244 64492 12284
rect 64012 11059 64052 11068
rect 64108 11864 64148 11873
rect 63915 11024 63957 11033
rect 63915 10984 63916 11024
rect 63956 10984 63957 11024
rect 63915 10975 63957 10984
rect 64108 11024 64148 11824
rect 64203 11864 64245 11873
rect 64203 11824 64204 11864
rect 64244 11824 64245 11864
rect 64203 11815 64245 11824
rect 64204 11192 64244 11815
rect 64300 11696 64340 12244
rect 64492 12235 64532 12244
rect 64395 12116 64437 12125
rect 64395 12076 64396 12116
rect 64436 12076 64437 12116
rect 64395 12067 64437 12076
rect 64300 11647 64340 11656
rect 64396 11696 64436 12067
rect 64588 11948 64628 11957
rect 64780 11948 64820 12496
rect 64628 11908 64820 11948
rect 64588 11899 64628 11908
rect 64876 11873 64916 14680
rect 65068 14671 65108 14680
rect 65163 14720 65205 14729
rect 65163 14680 65164 14720
rect 65204 14680 65205 14720
rect 65163 14671 65205 14680
rect 65356 14720 65396 14729
rect 65164 14586 65204 14671
rect 65068 14048 65108 14057
rect 65068 13376 65108 14008
rect 65164 13376 65204 13385
rect 65068 13336 65164 13376
rect 65164 13327 65204 13336
rect 65356 12980 65396 14680
rect 65931 14048 65973 14057
rect 65931 14008 65932 14048
rect 65972 14008 65973 14048
rect 65931 13999 65973 14008
rect 65932 13914 65972 13999
rect 65547 13880 65589 13889
rect 65547 13840 65548 13880
rect 65588 13840 65589 13880
rect 65547 13831 65589 13840
rect 65356 12940 65492 12980
rect 65164 12536 65204 12545
rect 64875 11864 64917 11873
rect 64875 11824 64876 11864
rect 64916 11824 64917 11864
rect 65164 11864 65204 12496
rect 65356 11864 65396 11873
rect 65164 11824 65356 11864
rect 64875 11815 64917 11824
rect 65356 11815 65396 11824
rect 65452 11789 65492 12940
rect 65548 12545 65588 13831
rect 65547 12536 65589 12545
rect 65547 12496 65548 12536
rect 65588 12496 65589 12536
rect 65547 12487 65589 12496
rect 66027 12536 66069 12545
rect 66027 12496 66028 12536
rect 66068 12496 66069 12536
rect 66027 12487 66069 12496
rect 64587 11780 64629 11789
rect 64587 11740 64588 11780
rect 64628 11740 64629 11780
rect 64587 11731 64629 11740
rect 64971 11780 65013 11789
rect 64971 11740 64972 11780
rect 65012 11740 65013 11780
rect 64971 11731 65013 11740
rect 65451 11780 65493 11789
rect 65451 11740 65452 11780
rect 65492 11740 65493 11780
rect 65451 11731 65493 11740
rect 64396 11647 64436 11656
rect 64588 11696 64628 11731
rect 64588 11645 64628 11656
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 64204 11152 64340 11192
rect 64108 10975 64148 10984
rect 63916 10890 63956 10975
rect 63820 10732 63956 10772
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 63435 10436 63477 10445
rect 63435 10396 63436 10436
rect 63476 10396 63477 10436
rect 63435 10387 63477 10396
rect 63436 10302 63476 10387
rect 63435 10184 63477 10193
rect 63435 10144 63436 10184
rect 63476 10144 63477 10184
rect 63435 10135 63477 10144
rect 63628 10184 63668 10195
rect 63436 10050 63476 10135
rect 63628 10109 63668 10144
rect 63724 10184 63764 10193
rect 63627 10100 63669 10109
rect 63627 10060 63628 10100
rect 63668 10060 63669 10100
rect 63627 10051 63669 10060
rect 63435 9512 63477 9521
rect 63435 9472 63436 9512
rect 63476 9472 63477 9512
rect 63435 9463 63477 9472
rect 63436 9378 63476 9463
rect 63724 9260 63764 10144
rect 63819 9260 63861 9269
rect 63724 9220 63820 9260
rect 63860 9220 63861 9260
rect 63819 9211 63861 9220
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 62859 8840 62901 8849
rect 62859 8800 62860 8840
rect 62900 8800 62901 8840
rect 62859 8791 62901 8800
rect 62860 8681 62900 8791
rect 62859 8672 62901 8681
rect 62859 8632 62860 8672
rect 62900 8632 62901 8672
rect 62859 8623 62901 8632
rect 63820 8672 63860 9211
rect 63820 8623 63860 8632
rect 63916 8672 63956 10732
rect 64203 10184 64245 10193
rect 64203 10144 64204 10184
rect 64244 10144 64245 10184
rect 64203 10135 64245 10144
rect 64300 10184 64340 11152
rect 64587 11024 64629 11033
rect 64587 10984 64588 11024
rect 64628 10984 64629 11024
rect 64587 10975 64629 10984
rect 64780 11024 64820 11033
rect 64588 10890 64628 10975
rect 64683 10940 64725 10949
rect 64683 10900 64684 10940
rect 64724 10900 64725 10940
rect 64683 10891 64725 10900
rect 64684 10772 64724 10891
rect 64587 10436 64629 10445
rect 64587 10396 64588 10436
rect 64628 10396 64629 10436
rect 64587 10387 64629 10396
rect 64300 10135 64340 10144
rect 64588 10184 64628 10387
rect 64684 10268 64724 10732
rect 64780 10436 64820 10984
rect 64972 11024 65012 11731
rect 64972 10975 65012 10984
rect 65164 11024 65204 11035
rect 65164 10949 65204 10984
rect 65260 11024 65300 11033
rect 65300 10984 65396 11024
rect 65260 10975 65300 10984
rect 65163 10940 65205 10949
rect 65163 10900 65164 10940
rect 65204 10900 65205 10940
rect 65163 10891 65205 10900
rect 64972 10772 65012 10781
rect 65012 10732 65300 10772
rect 64972 10723 65012 10732
rect 64972 10436 65012 10445
rect 64780 10396 64972 10436
rect 64972 10387 65012 10396
rect 64684 10228 65012 10268
rect 64588 10135 64628 10144
rect 64107 9008 64149 9017
rect 64107 8968 64108 9008
rect 64148 8968 64149 9008
rect 64107 8959 64149 8968
rect 63916 8623 63956 8632
rect 64011 8672 64053 8681
rect 64011 8632 64012 8672
rect 64052 8632 64053 8672
rect 64011 8623 64053 8632
rect 64108 8672 64148 8959
rect 64204 8672 64244 10135
rect 64684 10100 64724 10109
rect 64724 10060 64820 10100
rect 64684 10051 64724 10060
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 64588 9680 64628 9689
rect 64780 9680 64820 10060
rect 64628 9640 64820 9680
rect 64588 9631 64628 9640
rect 64875 9596 64917 9605
rect 64875 9556 64876 9596
rect 64916 9556 64917 9596
rect 64875 9547 64917 9556
rect 64780 9512 64820 9521
rect 64587 9260 64629 9269
rect 64587 9220 64588 9260
rect 64628 9220 64629 9260
rect 64587 9211 64629 9220
rect 64588 9126 64628 9211
rect 64780 9017 64820 9472
rect 64876 9462 64916 9547
rect 64972 9512 65012 10228
rect 65260 10184 65300 10732
rect 65260 10135 65300 10144
rect 65163 10100 65205 10109
rect 65163 10060 65164 10100
rect 65204 10060 65205 10100
rect 65163 10051 65205 10060
rect 64972 9463 65012 9472
rect 65068 9512 65108 9521
rect 64779 9008 64821 9017
rect 64779 8968 64780 9008
rect 64820 8968 64821 9008
rect 64779 8959 64821 8968
rect 65068 8849 65108 9472
rect 64395 8840 64437 8849
rect 64395 8800 64396 8840
rect 64436 8800 64437 8840
rect 64395 8791 64437 8800
rect 65067 8840 65109 8849
rect 65067 8800 65068 8840
rect 65108 8800 65109 8840
rect 65067 8791 65109 8800
rect 64300 8672 64340 8681
rect 64204 8632 64300 8672
rect 64108 8623 64148 8632
rect 64300 8623 64340 8632
rect 64012 8538 64052 8623
rect 64396 8588 64436 8791
rect 64780 8756 64820 8765
rect 64820 8716 65012 8756
rect 64780 8707 64820 8716
rect 64396 8539 64436 8548
rect 64492 8672 64532 8681
rect 64492 8513 64532 8632
rect 64588 8672 64628 8681
rect 64972 8672 65012 8716
rect 65164 8672 65204 10051
rect 65356 9596 65396 10984
rect 65451 10436 65493 10445
rect 65451 10396 65452 10436
rect 65492 10396 65493 10436
rect 65451 10387 65493 10396
rect 65356 9547 65396 9556
rect 65260 9512 65300 9521
rect 65260 9344 65300 9472
rect 65452 9512 65492 10387
rect 65452 9463 65492 9472
rect 65548 9344 65588 12487
rect 66028 11705 66068 12487
rect 66220 12041 66260 15427
rect 66508 14309 66548 16192
rect 66795 16183 66837 16192
rect 66892 16192 66988 16232
rect 66700 15560 66740 15569
rect 66507 14300 66549 14309
rect 66507 14260 66508 14300
rect 66548 14260 66549 14300
rect 66507 14251 66549 14260
rect 66700 14057 66740 15520
rect 66699 14048 66741 14057
rect 66699 14008 66700 14048
rect 66740 14008 66741 14048
rect 66699 13999 66741 14008
rect 66219 12032 66261 12041
rect 66219 11992 66220 12032
rect 66260 11992 66261 12032
rect 66219 11983 66261 11992
rect 66027 11696 66069 11705
rect 66027 11656 66028 11696
rect 66068 11656 66069 11696
rect 66027 11647 66069 11656
rect 65836 10856 65876 10865
rect 65644 10184 65684 10193
rect 65836 10184 65876 10816
rect 65684 10144 65876 10184
rect 66508 10184 66548 10193
rect 66548 10144 66644 10184
rect 65644 10135 65684 10144
rect 66508 10135 66548 10144
rect 66604 9521 66644 10144
rect 66796 9689 66836 16183
rect 66892 12629 66932 16192
rect 66988 16183 67028 16192
rect 67371 16232 67413 16241
rect 67371 16192 67372 16232
rect 67412 16192 67413 16232
rect 67371 16183 67413 16192
rect 67756 16232 67796 17116
rect 68055 17072 68095 17472
rect 68345 17156 68385 17472
rect 67852 17032 68095 17072
rect 68140 17116 68385 17156
rect 67852 16484 67892 17032
rect 67852 16435 67892 16444
rect 67275 16148 67317 16157
rect 67275 16108 67276 16148
rect 67316 16108 67317 16148
rect 67275 16099 67317 16108
rect 67179 14804 67221 14813
rect 67179 14764 67180 14804
rect 67220 14764 67221 14804
rect 67179 14755 67221 14764
rect 67180 14670 67220 14755
rect 67276 14552 67316 16099
rect 67372 16098 67412 16183
rect 67563 14636 67605 14645
rect 67563 14596 67564 14636
rect 67604 14596 67605 14636
rect 67563 14587 67605 14596
rect 67180 14512 67316 14552
rect 67372 14552 67412 14561
rect 67412 14512 67508 14552
rect 66987 14300 67029 14309
rect 66987 14260 66988 14300
rect 67028 14260 67029 14300
rect 66987 14251 67029 14260
rect 66891 12620 66933 12629
rect 66891 12580 66892 12620
rect 66932 12580 66933 12620
rect 66891 12571 66933 12580
rect 66891 10100 66933 10109
rect 66891 10060 66892 10100
rect 66932 10060 66933 10100
rect 66891 10051 66933 10060
rect 66795 9680 66837 9689
rect 66795 9640 66796 9680
rect 66836 9640 66837 9680
rect 66795 9631 66837 9640
rect 66892 9596 66932 10051
rect 66892 9547 66932 9556
rect 66603 9512 66645 9521
rect 66603 9472 66604 9512
rect 66644 9472 66645 9512
rect 66603 9463 66645 9472
rect 65260 9304 65588 9344
rect 66508 8840 66548 8849
rect 64972 8632 65204 8672
rect 66412 8800 66508 8840
rect 64491 8504 64533 8513
rect 64491 8464 64492 8504
rect 64532 8464 64533 8504
rect 64588 8504 64628 8632
rect 64875 8504 64917 8513
rect 64972 8504 65012 8513
rect 64588 8464 64820 8504
rect 64491 8455 64533 8464
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 62859 8168 62901 8177
rect 64108 8168 64148 8177
rect 62859 8128 62860 8168
rect 62900 8128 62901 8168
rect 62859 8119 62901 8128
rect 63628 8128 64108 8168
rect 62860 8034 62900 8119
rect 60940 7288 61076 7328
rect 61708 8000 61748 8009
rect 60843 7160 60885 7169
rect 60843 7120 60844 7160
rect 60884 7120 60885 7160
rect 60843 7111 60885 7120
rect 60748 7027 60788 7036
rect 60844 7026 60884 7111
rect 60651 6320 60693 6329
rect 60651 6280 60652 6320
rect 60692 6280 60693 6320
rect 60651 6271 60693 6280
rect 60940 6161 60980 7288
rect 61035 7160 61077 7169
rect 61035 7120 61036 7160
rect 61076 7120 61077 7160
rect 61035 7111 61077 7120
rect 61036 6488 61076 7111
rect 61324 6497 61364 6582
rect 61036 6439 61076 6448
rect 61228 6488 61268 6497
rect 61228 6320 61268 6448
rect 61323 6488 61365 6497
rect 61708 6488 61748 7960
rect 63628 8000 63668 8128
rect 64108 8119 64148 8128
rect 64780 8009 64820 8464
rect 64875 8464 64876 8504
rect 64916 8464 64972 8504
rect 64875 8455 64917 8464
rect 64972 8455 65012 8464
rect 63628 7951 63668 7960
rect 63819 8000 63861 8009
rect 63819 7960 63820 8000
rect 63860 7960 63861 8000
rect 63819 7951 63861 7960
rect 63916 8000 63956 8009
rect 63820 7866 63860 7951
rect 63052 7832 63092 7841
rect 62956 7792 63052 7832
rect 62187 7748 62229 7757
rect 62187 7708 62188 7748
rect 62228 7708 62229 7748
rect 62187 7699 62229 7708
rect 62188 7160 62228 7699
rect 62188 7111 62228 7120
rect 62572 7160 62612 7169
rect 62956 7160 62996 7792
rect 63052 7783 63092 7792
rect 63627 7748 63669 7757
rect 63627 7708 63628 7748
rect 63668 7708 63669 7748
rect 63627 7699 63669 7708
rect 63628 7614 63668 7699
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 62612 7120 62996 7160
rect 63436 7160 63476 7169
rect 63476 7120 63572 7160
rect 62572 7111 62612 7120
rect 63436 7111 63476 7120
rect 61323 6448 61324 6488
rect 61364 6448 61365 6488
rect 61323 6439 61365 6448
rect 61516 6448 61748 6488
rect 61899 6488 61941 6497
rect 61899 6448 61900 6488
rect 61940 6448 61941 6488
rect 61228 6280 61364 6320
rect 61036 6236 61076 6245
rect 61076 6196 61268 6236
rect 61036 6187 61076 6196
rect 60939 6152 60981 6161
rect 60939 6112 60940 6152
rect 60980 6112 60981 6152
rect 60939 6103 60981 6112
rect 61036 5816 61076 5825
rect 60651 5732 60693 5741
rect 60651 5692 60652 5732
rect 60692 5692 60693 5732
rect 60651 5683 60693 5692
rect 60404 5608 60500 5648
rect 60652 5648 60692 5683
rect 60171 5060 60213 5069
rect 60171 5020 60172 5060
rect 60212 5020 60213 5060
rect 60171 5011 60213 5020
rect 60075 4976 60117 4985
rect 60075 4936 60076 4976
rect 60116 4936 60117 4976
rect 60075 4927 60117 4936
rect 60076 4842 60116 4927
rect 60172 4304 60212 4313
rect 60076 4264 60172 4304
rect 59979 4220 60021 4229
rect 59979 4180 59980 4220
rect 60020 4180 60021 4220
rect 59979 4171 60021 4180
rect 59980 2969 60020 4171
rect 60076 3464 60116 4264
rect 60172 4255 60212 4264
rect 60076 3415 60116 3424
rect 60364 3053 60404 5608
rect 60652 5597 60692 5608
rect 60748 5564 60788 5573
rect 60459 5060 60501 5069
rect 60459 5020 60460 5060
rect 60500 5020 60501 5060
rect 60459 5011 60501 5020
rect 60363 3044 60405 3053
rect 60363 3004 60364 3044
rect 60404 3004 60405 3044
rect 60363 2995 60405 3004
rect 59979 2960 60021 2969
rect 59979 2920 59980 2960
rect 60020 2920 60021 2960
rect 59979 2911 60021 2920
rect 59980 1700 60020 2911
rect 60076 2792 60116 2801
rect 60076 2624 60116 2752
rect 60363 2708 60405 2717
rect 60363 2668 60364 2708
rect 60404 2668 60405 2708
rect 60363 2659 60405 2668
rect 60268 2624 60308 2633
rect 60076 2584 60268 2624
rect 60268 2575 60308 2584
rect 60364 2574 60404 2659
rect 60460 2624 60500 5011
rect 60748 4145 60788 5524
rect 61036 5153 61076 5776
rect 61228 5648 61268 6196
rect 61324 5657 61364 6280
rect 61516 5657 61556 6448
rect 61899 6439 61941 6448
rect 61708 6320 61748 6329
rect 61228 5599 61268 5608
rect 61323 5648 61365 5657
rect 61323 5608 61324 5648
rect 61364 5608 61365 5648
rect 61323 5599 61365 5608
rect 61515 5648 61557 5657
rect 61515 5608 61516 5648
rect 61556 5608 61557 5648
rect 61515 5599 61557 5608
rect 61612 5648 61652 5657
rect 61708 5648 61748 6280
rect 61652 5608 61748 5648
rect 61612 5599 61652 5608
rect 61035 5144 61077 5153
rect 61035 5104 61036 5144
rect 61076 5104 61077 5144
rect 61035 5095 61077 5104
rect 60939 4976 60981 4985
rect 60939 4936 60940 4976
rect 60980 4936 60981 4976
rect 60939 4927 60981 4936
rect 60747 4136 60789 4145
rect 60747 4096 60748 4136
rect 60788 4096 60789 4136
rect 60747 4087 60789 4096
rect 60940 3464 60980 4927
rect 61324 4808 61364 5599
rect 61419 5144 61461 5153
rect 61419 5104 61420 5144
rect 61460 5104 61461 5144
rect 61419 5095 61461 5104
rect 61420 4976 61460 5095
rect 61516 4985 61556 5599
rect 61611 5060 61653 5069
rect 61611 5020 61612 5060
rect 61652 5020 61653 5060
rect 61611 5011 61653 5020
rect 61900 5060 61940 6439
rect 63436 6320 63476 6331
rect 63436 6245 63476 6280
rect 63435 6236 63477 6245
rect 63435 6196 63436 6236
rect 63476 6196 63477 6236
rect 63435 6187 63477 6196
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 63339 5900 63381 5909
rect 63339 5860 63340 5900
rect 63380 5860 63381 5900
rect 63339 5851 63381 5860
rect 61995 5732 62037 5741
rect 61995 5692 61996 5732
rect 62036 5692 62037 5732
rect 61995 5683 62037 5692
rect 61900 5011 61940 5020
rect 61420 4927 61460 4936
rect 61515 4976 61557 4985
rect 61515 4936 61516 4976
rect 61556 4936 61557 4976
rect 61515 4927 61557 4936
rect 61612 4976 61652 5011
rect 61612 4901 61652 4936
rect 61804 4976 61844 4985
rect 61611 4892 61653 4901
rect 61611 4852 61612 4892
rect 61652 4852 61653 4892
rect 61611 4843 61653 4852
rect 61516 4808 61556 4817
rect 61612 4812 61652 4843
rect 61324 4768 61516 4808
rect 61516 4759 61556 4768
rect 61228 4724 61268 4733
rect 61228 4145 61268 4684
rect 61804 4313 61844 4936
rect 61996 4976 62036 5683
rect 62475 5648 62517 5657
rect 62475 5608 62476 5648
rect 62516 5608 62517 5648
rect 62475 5599 62517 5608
rect 62476 5514 62516 5599
rect 62955 5480 62997 5489
rect 62955 5440 62956 5480
rect 62996 5440 62997 5480
rect 62955 5431 62997 5440
rect 62956 5060 62996 5431
rect 62956 5011 62996 5020
rect 61996 4927 62036 4936
rect 63340 4976 63380 5851
rect 63532 5657 63572 7120
rect 63916 7085 63956 7960
rect 64204 8000 64244 8009
rect 64107 7160 64149 7169
rect 64107 7120 64108 7160
rect 64148 7120 64149 7160
rect 64107 7111 64149 7120
rect 63915 7076 63957 7085
rect 63915 7036 63916 7076
rect 63956 7036 63957 7076
rect 63915 7027 63957 7036
rect 63915 6740 63957 6749
rect 63915 6700 63916 6740
rect 63956 6700 63957 6740
rect 63915 6691 63957 6700
rect 63627 5732 63669 5741
rect 63627 5692 63628 5732
rect 63668 5692 63669 5732
rect 63627 5683 63669 5692
rect 63531 5648 63573 5657
rect 63531 5608 63532 5648
rect 63572 5608 63573 5648
rect 63531 5599 63573 5608
rect 63628 5573 63668 5683
rect 63627 5564 63669 5573
rect 63627 5524 63628 5564
rect 63668 5524 63669 5564
rect 63627 5515 63669 5524
rect 63628 5480 63668 5515
rect 63628 5429 63668 5440
rect 63916 4985 63956 6691
rect 64108 6497 64148 7111
rect 64107 6488 64149 6497
rect 64107 6448 64108 6488
rect 64148 6448 64149 6488
rect 64107 6439 64149 6448
rect 64204 5825 64244 7960
rect 64300 8000 64340 8009
rect 64300 7169 64340 7960
rect 64395 8000 64437 8009
rect 64395 7960 64396 8000
rect 64436 7960 64437 8000
rect 64395 7951 64437 7960
rect 64684 8000 64724 8009
rect 64396 7412 64436 7951
rect 64684 7841 64724 7960
rect 64779 8000 64821 8009
rect 64779 7960 64780 8000
rect 64820 7960 64821 8000
rect 64779 7951 64821 7960
rect 64683 7832 64725 7841
rect 64683 7792 64684 7832
rect 64724 7792 64725 7832
rect 64876 7832 64916 8455
rect 65644 8168 65684 8177
rect 64972 8128 65204 8168
rect 64972 8000 65012 8128
rect 64972 7951 65012 7960
rect 65067 8000 65109 8009
rect 65067 7960 65068 8000
rect 65108 7960 65109 8000
rect 65067 7951 65109 7960
rect 65068 7866 65108 7951
rect 64876 7792 65012 7832
rect 64683 7783 64725 7792
rect 64588 7412 64628 7421
rect 64396 7372 64588 7412
rect 64588 7363 64628 7372
rect 64972 7169 65012 7792
rect 65164 7757 65204 8128
rect 65684 8128 65972 8168
rect 65644 8119 65684 8128
rect 65932 8084 65972 8128
rect 66028 8084 66068 8093
rect 65932 8044 66028 8084
rect 66028 8035 66068 8044
rect 65547 8000 65589 8009
rect 65547 7960 65548 8000
rect 65588 7960 65589 8000
rect 65547 7951 65589 7960
rect 65740 8000 65780 8011
rect 65259 7916 65301 7925
rect 65259 7876 65260 7916
rect 65300 7876 65301 7916
rect 65259 7867 65301 7876
rect 65163 7748 65205 7757
rect 65163 7708 65164 7748
rect 65204 7708 65205 7748
rect 65163 7699 65205 7708
rect 65260 7412 65300 7867
rect 65548 7866 65588 7951
rect 65740 7925 65780 7960
rect 65836 8000 65876 8009
rect 65739 7916 65781 7925
rect 65739 7876 65740 7916
rect 65780 7876 65781 7916
rect 65739 7867 65781 7876
rect 65643 7832 65685 7841
rect 65643 7792 65644 7832
rect 65684 7792 65685 7832
rect 65643 7783 65685 7792
rect 65356 7748 65396 7757
rect 65396 7708 65492 7748
rect 65356 7699 65396 7708
rect 65356 7412 65396 7421
rect 65260 7372 65356 7412
rect 65356 7363 65396 7372
rect 64299 7160 64341 7169
rect 64299 7120 64300 7160
rect 64340 7120 64341 7160
rect 64299 7111 64341 7120
rect 64780 7160 64820 7169
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 64780 6749 64820 7120
rect 64971 7160 65013 7169
rect 64971 7120 64972 7160
rect 65012 7120 65013 7160
rect 64971 7111 65013 7120
rect 65068 7160 65108 7169
rect 65260 7160 65300 7169
rect 65108 7120 65204 7160
rect 65068 7111 65108 7120
rect 64875 7076 64917 7085
rect 64875 7036 64876 7076
rect 64916 7036 64917 7076
rect 64875 7027 64917 7036
rect 64876 6942 64916 7027
rect 64972 7026 65012 7111
rect 64779 6740 64821 6749
rect 64779 6700 64780 6740
rect 64820 6700 64821 6740
rect 64779 6691 64821 6700
rect 65164 6656 65204 7120
rect 65260 6917 65300 7120
rect 65452 7160 65492 7708
rect 65452 7111 65492 7120
rect 65259 6908 65301 6917
rect 65259 6868 65260 6908
rect 65300 6868 65301 6908
rect 65259 6859 65301 6868
rect 65547 6908 65589 6917
rect 65547 6868 65548 6908
rect 65588 6868 65589 6908
rect 65547 6859 65589 6868
rect 65164 6616 65396 6656
rect 65259 6488 65301 6497
rect 65259 6448 65260 6488
rect 65300 6448 65301 6488
rect 65259 6439 65301 6448
rect 64203 5816 64245 5825
rect 64012 5776 64204 5816
rect 64244 5776 64245 5816
rect 63340 4927 63380 4936
rect 63627 4976 63669 4985
rect 63627 4936 63628 4976
rect 63668 4936 63669 4976
rect 63627 4927 63669 4936
rect 63915 4976 63957 4985
rect 63915 4936 63916 4976
rect 63956 4936 63957 4976
rect 63915 4927 63957 4936
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 61803 4304 61845 4313
rect 61803 4264 61804 4304
rect 61844 4264 61845 4304
rect 61803 4255 61845 4264
rect 62763 4304 62805 4313
rect 62763 4264 62764 4304
rect 62804 4264 62805 4304
rect 62763 4255 62805 4264
rect 61227 4136 61269 4145
rect 61227 4096 61228 4136
rect 61268 4096 61269 4136
rect 61227 4087 61269 4096
rect 60555 3128 60597 3137
rect 60555 3088 60556 3128
rect 60596 3088 60597 3128
rect 60555 3079 60597 3088
rect 60460 2575 60500 2584
rect 60459 1952 60501 1961
rect 60459 1912 60460 1952
rect 60500 1912 60501 1952
rect 60459 1903 60501 1912
rect 60460 1818 60500 1903
rect 59980 1660 60500 1700
rect 59116 1063 59156 1072
rect 59883 1112 59925 1121
rect 59883 1072 59884 1112
rect 59924 1072 59925 1112
rect 59883 1063 59925 1072
rect 60075 1112 60117 1121
rect 60075 1072 60076 1112
rect 60116 1072 60117 1112
rect 60075 1063 60117 1072
rect 60460 1112 60500 1660
rect 60556 1205 60596 3079
rect 60651 2540 60693 2549
rect 60651 2500 60652 2540
rect 60692 2500 60693 2540
rect 60651 2491 60693 2500
rect 60555 1196 60597 1205
rect 60555 1156 60556 1196
rect 60596 1156 60597 1196
rect 60555 1147 60597 1156
rect 60460 1063 60500 1072
rect 60556 1112 60596 1147
rect 60076 978 60116 1063
rect 60556 1062 60596 1072
rect 60652 1112 60692 2491
rect 60940 1961 60980 3424
rect 61804 2900 61844 4255
rect 62091 3716 62133 3725
rect 62091 3676 62092 3716
rect 62132 3676 62133 3716
rect 62091 3667 62133 3676
rect 62092 3632 62132 3667
rect 62092 3581 62132 3592
rect 62764 2969 62804 4255
rect 63244 4136 63284 4145
rect 62860 4052 62900 4061
rect 62860 3641 62900 4012
rect 63244 3716 63284 4096
rect 63244 3676 63380 3716
rect 62859 3632 62901 3641
rect 62859 3592 62860 3632
rect 62900 3592 62901 3632
rect 62859 3583 62901 3592
rect 63340 3338 63380 3676
rect 63340 3289 63380 3298
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 62763 2960 62805 2969
rect 62763 2920 62764 2960
rect 62804 2920 62805 2960
rect 62763 2911 62805 2920
rect 61804 2860 61940 2900
rect 61611 2540 61653 2549
rect 61611 2500 61612 2540
rect 61652 2500 61653 2540
rect 61611 2491 61653 2500
rect 61612 2120 61652 2491
rect 61612 2071 61652 2080
rect 60939 1952 60981 1961
rect 60939 1912 60940 1952
rect 60980 1912 60981 1952
rect 60939 1903 60981 1912
rect 61804 1952 61844 1961
rect 61612 1700 61652 1709
rect 60843 1280 60885 1289
rect 60843 1240 60844 1280
rect 60884 1240 60885 1280
rect 60843 1231 60885 1240
rect 60844 1146 60884 1231
rect 61612 1112 61652 1660
rect 61804 1373 61844 1912
rect 61803 1364 61845 1373
rect 61803 1324 61804 1364
rect 61844 1324 61845 1364
rect 61803 1315 61845 1324
rect 61708 1112 61748 1121
rect 61612 1072 61708 1112
rect 60652 1063 60692 1072
rect 61708 1063 61748 1072
rect 61804 1112 61844 1121
rect 61900 1112 61940 2860
rect 62188 2792 62228 2801
rect 62188 1952 62228 2752
rect 62188 1903 62228 1912
rect 62475 1364 62517 1373
rect 62475 1324 62476 1364
rect 62516 1324 62517 1364
rect 62475 1315 62517 1324
rect 61996 1280 62036 1289
rect 62283 1280 62325 1289
rect 62036 1240 62228 1280
rect 61996 1231 62036 1240
rect 61844 1072 61940 1112
rect 61996 1112 62036 1123
rect 61804 1063 61844 1072
rect 61996 1037 62036 1072
rect 62188 1112 62228 1240
rect 62283 1240 62284 1280
rect 62324 1240 62325 1280
rect 62283 1231 62325 1240
rect 62188 1063 62228 1072
rect 62284 1112 62324 1231
rect 62476 1230 62516 1315
rect 62284 1063 62324 1072
rect 62476 1112 62516 1121
rect 62668 1112 62708 1121
rect 62516 1072 62668 1112
rect 62476 1063 62516 1072
rect 62668 1063 62708 1072
rect 62764 1112 62804 2911
rect 63628 2900 63668 4927
rect 64012 4313 64052 5776
rect 64203 5767 64245 5776
rect 64587 5816 64629 5825
rect 64587 5776 64588 5816
rect 64628 5776 64629 5816
rect 64587 5767 64629 5776
rect 65067 5816 65109 5825
rect 65067 5776 65068 5816
rect 65108 5776 65109 5816
rect 65067 5767 65109 5776
rect 64203 5648 64245 5657
rect 64203 5608 64204 5648
rect 64244 5608 64245 5648
rect 64203 5599 64245 5608
rect 64588 5648 64628 5767
rect 64588 5599 64628 5608
rect 64779 5648 64821 5657
rect 64779 5608 64780 5648
rect 64820 5608 64821 5648
rect 64779 5599 64821 5608
rect 64876 5648 64916 5657
rect 64204 4976 64244 5599
rect 64684 5489 64724 5574
rect 64780 5514 64820 5599
rect 64683 5480 64725 5489
rect 64683 5440 64684 5480
rect 64724 5440 64725 5480
rect 64683 5431 64725 5440
rect 64779 5396 64821 5405
rect 64779 5356 64780 5396
rect 64820 5356 64821 5396
rect 64779 5347 64821 5356
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 64011 4304 64053 4313
rect 64011 4264 64012 4304
rect 64052 4264 64053 4304
rect 64011 4255 64053 4264
rect 64012 3800 64052 4255
rect 64108 4136 64148 4145
rect 64204 4136 64244 4936
rect 64148 4096 64244 4136
rect 64108 4087 64148 4096
rect 64352 3800 64720 3809
rect 64012 3760 64244 3800
rect 64011 3632 64053 3641
rect 64011 3592 64012 3632
rect 64052 3592 64053 3632
rect 64204 3632 64244 3760
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 64780 3632 64820 5347
rect 64876 5153 64916 5608
rect 65068 5648 65108 5767
rect 65163 5732 65205 5741
rect 65163 5692 65164 5732
rect 65204 5692 65205 5732
rect 65163 5683 65205 5692
rect 65068 5599 65108 5608
rect 65164 5648 65204 5683
rect 65164 5597 65204 5608
rect 65260 5648 65300 6439
rect 65356 6329 65396 6616
rect 65355 6320 65397 6329
rect 65355 6280 65356 6320
rect 65396 6280 65397 6320
rect 65355 6271 65397 6280
rect 65260 5405 65300 5608
rect 65356 5648 65396 6271
rect 65259 5396 65301 5405
rect 65259 5356 65260 5396
rect 65300 5356 65301 5396
rect 65259 5347 65301 5356
rect 64875 5144 64917 5153
rect 64875 5104 64876 5144
rect 64916 5104 64917 5144
rect 64875 5095 64917 5104
rect 65356 5144 65396 5608
rect 65548 5489 65588 6859
rect 65644 6488 65684 7783
rect 65836 7412 65876 7960
rect 66412 8000 66452 8800
rect 66508 8791 66548 8800
rect 66604 8681 66644 9463
rect 66603 8672 66645 8681
rect 66603 8632 66604 8672
rect 66644 8632 66645 8672
rect 66603 8623 66645 8632
rect 66412 7951 66452 7960
rect 66988 7916 67028 14251
rect 67083 13964 67125 13973
rect 67083 13924 67084 13964
rect 67124 13924 67125 13964
rect 67083 13915 67125 13924
rect 67084 13830 67124 13915
rect 67180 12980 67220 14512
rect 67372 14503 67412 14512
rect 67276 14048 67316 14059
rect 67276 13973 67316 14008
rect 67372 14048 67412 14057
rect 67275 13964 67317 13973
rect 67275 13924 67276 13964
rect 67316 13924 67317 13964
rect 67275 13915 67317 13924
rect 67372 13889 67412 14008
rect 67468 14048 67508 14512
rect 67564 14502 67604 14587
rect 67564 14048 67604 14057
rect 67468 14008 67564 14048
rect 67371 13880 67413 13889
rect 67371 13840 67372 13880
rect 67412 13840 67413 13880
rect 67371 13831 67413 13840
rect 67468 13301 67508 14008
rect 67564 13999 67604 14008
rect 67563 13880 67605 13889
rect 67563 13840 67564 13880
rect 67604 13840 67605 13880
rect 67563 13831 67605 13840
rect 67564 13746 67604 13831
rect 67467 13292 67509 13301
rect 67467 13252 67468 13292
rect 67508 13252 67509 13292
rect 67467 13243 67509 13252
rect 67756 12980 67796 16192
rect 67947 16232 67989 16241
rect 67947 16192 67948 16232
rect 67988 16192 67989 16232
rect 67947 16183 67989 16192
rect 68140 16232 68180 17116
rect 68455 17072 68495 17472
rect 68745 17156 68785 17472
rect 68236 17032 68495 17072
rect 68716 17116 68785 17156
rect 68236 16484 68276 17032
rect 68236 16435 68276 16444
rect 67851 15728 67893 15737
rect 67851 15688 67852 15728
rect 67892 15688 67893 15728
rect 67851 15679 67893 15688
rect 67852 15594 67892 15679
rect 67948 15476 67988 16183
rect 67852 15436 67988 15476
rect 67852 13721 67892 15436
rect 68044 15392 68084 15401
rect 67948 14720 67988 14729
rect 68044 14720 68084 15352
rect 67988 14680 68084 14720
rect 67948 14671 67988 14680
rect 68140 14552 68180 16192
rect 68524 16232 68564 16241
rect 68716 16232 68756 17116
rect 68855 17072 68895 17472
rect 69145 17156 69185 17472
rect 68564 16192 68756 16232
rect 68812 17032 68895 17072
rect 69004 17116 69185 17156
rect 68524 16073 68564 16192
rect 68523 16064 68565 16073
rect 68523 16024 68524 16064
rect 68564 16024 68565 16064
rect 68523 16015 68565 16024
rect 68620 16064 68660 16073
rect 68812 16064 68852 17032
rect 69004 16241 69044 17116
rect 69255 17072 69295 17472
rect 69545 17156 69585 17472
rect 69100 17032 69295 17072
rect 69388 17116 69585 17156
rect 69100 16484 69140 17032
rect 69100 16435 69140 16444
rect 69003 16232 69045 16241
rect 69003 16192 69004 16232
rect 69044 16192 69045 16232
rect 69003 16183 69045 16192
rect 69388 16232 69428 17116
rect 69655 17072 69695 17472
rect 69945 17156 69985 17472
rect 69484 17032 69695 17072
rect 69772 17116 69985 17156
rect 69484 16484 69524 17032
rect 69484 16435 69524 16444
rect 69004 16098 69044 16183
rect 69388 16157 69428 16192
rect 69772 16232 69812 17116
rect 70055 17072 70095 17472
rect 70345 17240 70385 17472
rect 69868 17032 70095 17072
rect 70156 17200 70385 17240
rect 69868 16484 69908 17032
rect 69868 16435 69908 16444
rect 70156 16241 70196 17200
rect 70455 17072 70495 17472
rect 70745 17156 70785 17472
rect 70252 17032 70495 17072
rect 70540 17116 70785 17156
rect 70252 16484 70292 17032
rect 70540 16988 70580 17116
rect 70855 17072 70895 17472
rect 71145 17156 71185 17472
rect 70444 16948 70580 16988
rect 70636 17032 70895 17072
rect 70937 17116 71185 17156
rect 70444 16652 70484 16948
rect 70444 16612 70567 16652
rect 70252 16435 70292 16444
rect 69387 16148 69429 16157
rect 69387 16108 69388 16148
rect 69428 16108 69429 16148
rect 69387 16099 69429 16108
rect 68660 16024 68852 16064
rect 68620 16015 68660 16024
rect 69772 15989 69812 16192
rect 70155 16232 70197 16241
rect 70155 16192 70156 16232
rect 70196 16192 70197 16232
rect 70155 16183 70197 16192
rect 70527 16221 70567 16612
rect 70636 16484 70676 17032
rect 70937 16988 70977 17116
rect 71255 17072 71295 17472
rect 71403 17156 71445 17165
rect 71545 17156 71585 17472
rect 71655 17165 71695 17472
rect 71403 17116 71404 17156
rect 71444 17116 71445 17156
rect 71403 17107 71445 17116
rect 71500 17116 71585 17156
rect 71654 17156 71696 17165
rect 71945 17156 71985 17472
rect 71654 17116 71655 17156
rect 71695 17116 71696 17156
rect 70636 16435 70676 16444
rect 70924 16948 70977 16988
rect 71020 17032 71295 17072
rect 70156 16098 70196 16183
rect 70527 16073 70567 16181
rect 70924 16232 70964 16948
rect 71020 16484 71060 17032
rect 71020 16435 71060 16444
rect 71404 16484 71444 17107
rect 71404 16435 71444 16444
rect 70526 16064 70568 16073
rect 70526 16024 70527 16064
rect 70567 16024 70568 16064
rect 70526 16015 70568 16024
rect 69099 15980 69141 15989
rect 69099 15940 69100 15980
rect 69140 15940 69141 15980
rect 69099 15931 69141 15940
rect 69771 15980 69813 15989
rect 69771 15940 69772 15980
rect 69812 15940 69813 15980
rect 69771 15931 69813 15940
rect 68715 15476 68757 15485
rect 68715 15436 68716 15476
rect 68756 15436 68757 15476
rect 68715 15427 68757 15436
rect 68716 15342 68756 15427
rect 68908 15308 68948 15317
rect 68908 14888 68948 15268
rect 68716 14848 68948 14888
rect 68235 14636 68277 14645
rect 68235 14596 68236 14636
rect 68276 14596 68277 14636
rect 68235 14587 68277 14596
rect 67948 14512 68180 14552
rect 67851 13712 67893 13721
rect 67851 13672 67852 13712
rect 67892 13672 67893 13712
rect 67851 13663 67893 13672
rect 67180 12940 67316 12980
rect 67756 12940 67892 12980
rect 67179 12788 67221 12797
rect 67179 12748 67180 12788
rect 67220 12748 67221 12788
rect 67179 12739 67221 12748
rect 67180 12704 67220 12739
rect 67180 12461 67220 12664
rect 67179 12452 67221 12461
rect 67179 12412 67180 12452
rect 67220 12412 67221 12452
rect 67179 12403 67221 12412
rect 67276 10520 67316 12940
rect 67372 12536 67412 12545
rect 67756 12536 67796 12545
rect 67372 11621 67412 12496
rect 67564 12496 67756 12536
rect 67564 11864 67604 12496
rect 67756 12487 67796 12496
rect 67564 11815 67604 11824
rect 67371 11612 67413 11621
rect 67371 11572 67372 11612
rect 67412 11572 67413 11612
rect 67371 11563 67413 11572
rect 67852 10520 67892 12940
rect 67276 10480 67412 10520
rect 67275 10352 67317 10361
rect 67275 10312 67276 10352
rect 67316 10312 67317 10352
rect 67275 10303 67317 10312
rect 67276 9512 67316 10303
rect 67276 9463 67316 9472
rect 67275 8672 67317 8681
rect 67275 8632 67276 8672
rect 67316 8632 67317 8672
rect 67275 8623 67317 8632
rect 67276 8000 67316 8623
rect 67276 7951 67316 7960
rect 66892 7876 67028 7916
rect 66027 7748 66069 7757
rect 66027 7708 66028 7748
rect 66068 7708 66069 7748
rect 66027 7699 66069 7708
rect 65932 7412 65972 7421
rect 65836 7372 65932 7412
rect 65932 7363 65972 7372
rect 65836 7169 65876 7255
rect 65739 7160 65781 7169
rect 65739 7120 65740 7160
rect 65780 7120 65781 7160
rect 65739 7111 65781 7120
rect 65835 7161 65877 7169
rect 65835 7120 65836 7161
rect 65876 7120 65877 7161
rect 65835 7111 65877 7120
rect 66028 7160 66068 7699
rect 66028 7111 66068 7120
rect 66220 7160 66260 7169
rect 65547 5480 65589 5489
rect 65547 5440 65548 5480
rect 65588 5440 65589 5480
rect 65547 5431 65589 5440
rect 65644 5312 65684 6448
rect 65356 5095 65396 5104
rect 65452 5272 65684 5312
rect 65163 5060 65205 5069
rect 65163 5020 65164 5060
rect 65204 5020 65205 5060
rect 65163 5011 65205 5020
rect 64204 3592 64436 3632
rect 64011 3583 64053 3592
rect 64012 3498 64052 3583
rect 63820 3464 63860 3473
rect 63820 2900 63860 3424
rect 63915 3464 63957 3473
rect 63915 3424 63916 3464
rect 63956 3424 63957 3464
rect 63915 3415 63957 3424
rect 64108 3464 64148 3473
rect 64300 3464 64340 3473
rect 64148 3424 64300 3464
rect 64108 3415 64148 3424
rect 64300 3415 64340 3424
rect 64396 3464 64436 3592
rect 64396 3415 64436 3424
rect 64492 3592 64820 3632
rect 64492 3464 64532 3592
rect 64492 3415 64532 3424
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 63916 3330 63956 3415
rect 64588 3330 64628 3415
rect 64107 3296 64149 3305
rect 64107 3256 64108 3296
rect 64148 3256 64149 3296
rect 64107 3247 64149 3256
rect 63628 2860 63764 2900
rect 63820 2876 64052 2900
rect 63820 2860 64012 2876
rect 63051 1952 63093 1961
rect 63051 1912 63052 1952
rect 63092 1912 63093 1952
rect 63051 1903 63093 1912
rect 63052 1818 63092 1903
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 62859 1196 62901 1205
rect 62859 1156 62860 1196
rect 62900 1156 62901 1196
rect 62859 1147 62901 1156
rect 62764 1063 62804 1072
rect 62860 1112 62900 1147
rect 62860 1061 62900 1072
rect 62956 1112 62996 1121
rect 61995 1028 62037 1037
rect 61995 988 61996 1028
rect 62036 988 62037 1028
rect 61995 979 62037 988
rect 62956 953 62996 1072
rect 63628 1037 63668 2860
rect 63724 2792 63764 2860
rect 64012 2796 64052 2836
rect 63724 2752 63956 2792
rect 63724 2624 63764 2633
rect 63627 1028 63669 1037
rect 63627 988 63628 1028
rect 63668 988 63669 1028
rect 63627 979 63669 988
rect 63724 953 63764 2584
rect 63820 2624 63860 2633
rect 63916 2624 63956 2752
rect 64012 2624 64052 2633
rect 63916 2584 64012 2624
rect 63820 2465 63860 2584
rect 64012 2575 64052 2584
rect 63819 2456 63861 2465
rect 63819 2416 63820 2456
rect 63860 2416 63861 2456
rect 63819 2407 63861 2416
rect 64108 2036 64148 3247
rect 65164 2900 65204 5011
rect 65452 4136 65492 5272
rect 65643 5144 65685 5153
rect 65643 5104 65644 5144
rect 65684 5104 65685 5144
rect 65643 5095 65685 5104
rect 65644 5010 65684 5095
rect 65740 4985 65780 7111
rect 66220 6917 66260 7120
rect 66412 7160 66452 7169
rect 66316 7076 66356 7085
rect 66219 6908 66261 6917
rect 66219 6868 66220 6908
rect 66260 6868 66261 6908
rect 66219 6859 66261 6868
rect 65836 6616 66068 6656
rect 65836 6329 65876 6616
rect 66028 6572 66068 6616
rect 66028 6523 66068 6532
rect 65931 6488 65973 6497
rect 66316 6488 66356 7036
rect 65931 6448 65932 6488
rect 65972 6448 65973 6488
rect 65931 6439 65973 6448
rect 66220 6448 66356 6488
rect 65932 6354 65972 6439
rect 65835 6320 65877 6329
rect 65835 6280 65836 6320
rect 65876 6280 65877 6320
rect 65835 6271 65877 6280
rect 66220 5657 66260 6448
rect 66316 6320 66356 6329
rect 66412 6320 66452 7120
rect 66603 7160 66645 7169
rect 66603 7120 66604 7160
rect 66644 7120 66645 7160
rect 66603 7111 66645 7120
rect 66796 7160 66836 7171
rect 66604 7026 66644 7111
rect 66796 7085 66836 7120
rect 66700 7076 66740 7085
rect 66356 6280 66452 6320
rect 66604 6488 66644 6497
rect 66316 6271 66356 6280
rect 66316 5900 66356 5909
rect 66604 5900 66644 6448
rect 66356 5860 66644 5900
rect 66316 5851 66356 5860
rect 66219 5648 66261 5657
rect 66219 5608 66220 5648
rect 66260 5608 66261 5648
rect 66507 5648 66549 5657
rect 66219 5599 66261 5608
rect 66316 5606 66356 5615
rect 66507 5608 66508 5648
rect 66548 5608 66549 5648
rect 66507 5599 66549 5608
rect 66604 5648 66644 5657
rect 66700 5648 66740 7036
rect 66795 7076 66837 7085
rect 66795 7036 66796 7076
rect 66836 7036 66837 7076
rect 66795 7027 66837 7036
rect 66796 6497 66836 7027
rect 66795 6488 66837 6497
rect 66795 6448 66796 6488
rect 66836 6448 66837 6488
rect 66795 6439 66837 6448
rect 66644 5608 66740 5648
rect 66604 5599 66644 5608
rect 66316 5489 66356 5566
rect 66508 5514 66548 5599
rect 66123 5480 66165 5489
rect 66123 5440 66124 5480
rect 66164 5440 66165 5480
rect 66123 5431 66165 5440
rect 66315 5480 66357 5489
rect 66315 5440 66316 5480
rect 66356 5440 66357 5480
rect 66315 5431 66357 5440
rect 66124 5069 66164 5431
rect 66316 5144 66356 5431
rect 66316 5104 66452 5144
rect 66123 5060 66165 5069
rect 66123 5020 66124 5060
rect 66164 5020 66165 5060
rect 66123 5011 66165 5020
rect 65547 4976 65589 4985
rect 65547 4936 65548 4976
rect 65588 4936 65589 4976
rect 65547 4927 65589 4936
rect 65739 4976 65781 4985
rect 65739 4936 65740 4976
rect 65780 4936 65781 4976
rect 65739 4927 65781 4936
rect 65836 4976 65876 4985
rect 66124 4976 66164 5011
rect 65876 4936 65972 4976
rect 65836 4927 65876 4936
rect 65548 4842 65588 4927
rect 65548 4136 65588 4145
rect 65452 4096 65548 4136
rect 65260 4061 65300 4092
rect 65259 4052 65301 4061
rect 65259 4012 65260 4052
rect 65300 4012 65301 4052
rect 65259 4003 65301 4012
rect 65260 3968 65300 4003
rect 65260 3473 65300 3928
rect 65259 3464 65301 3473
rect 65259 3424 65260 3464
rect 65300 3424 65301 3464
rect 65259 3415 65301 3424
rect 65452 3305 65492 4096
rect 65548 4087 65588 4096
rect 65451 3296 65493 3305
rect 65451 3256 65452 3296
rect 65492 3256 65493 3296
rect 65451 3247 65493 3256
rect 64203 2876 64245 2885
rect 64203 2836 64204 2876
rect 64244 2836 64245 2876
rect 65164 2860 65300 2900
rect 64203 2827 64245 2836
rect 64204 2624 64244 2827
rect 64780 2717 64820 2802
rect 64491 2708 64533 2717
rect 64491 2668 64492 2708
rect 64532 2668 64533 2708
rect 64491 2659 64533 2668
rect 64779 2708 64821 2717
rect 64779 2668 64780 2708
rect 64820 2668 64821 2708
rect 64779 2659 64821 2668
rect 64204 2575 64244 2584
rect 64396 2624 64436 2635
rect 64396 2549 64436 2584
rect 64492 2624 64532 2659
rect 64492 2573 64532 2584
rect 64684 2624 64724 2633
rect 64395 2540 64437 2549
rect 64395 2500 64396 2540
rect 64436 2500 64437 2540
rect 64395 2491 64437 2500
rect 64684 2465 64724 2584
rect 64876 2624 64916 2633
rect 64916 2584 65204 2624
rect 64876 2575 64916 2584
rect 64779 2540 64821 2549
rect 64779 2500 64780 2540
rect 64820 2500 64821 2540
rect 64779 2491 64821 2500
rect 64300 2456 64340 2465
rect 64204 2416 64300 2456
rect 64204 2120 64244 2416
rect 64300 2407 64340 2416
rect 64683 2456 64725 2465
rect 64683 2416 64684 2456
rect 64724 2416 64725 2456
rect 64683 2407 64725 2416
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 64204 2080 64532 2120
rect 64012 1996 64148 2036
rect 64492 2036 64532 2080
rect 63820 1112 63860 1121
rect 64012 1112 64052 1996
rect 64492 1987 64532 1996
rect 64204 1700 64244 1709
rect 64107 1448 64149 1457
rect 64107 1408 64108 1448
rect 64148 1408 64149 1448
rect 64107 1399 64149 1408
rect 63860 1072 64052 1112
rect 64108 1112 64148 1399
rect 63820 1063 63860 1072
rect 64108 1063 64148 1072
rect 64204 1028 64244 1660
rect 64780 1289 64820 2491
rect 65164 2129 65204 2584
rect 65163 2120 65205 2129
rect 65163 2080 65164 2120
rect 65204 2080 65205 2120
rect 65163 2071 65205 2080
rect 64876 1952 64916 1961
rect 64916 1912 65108 1952
rect 64876 1903 64916 1912
rect 64492 1280 64532 1289
rect 64779 1280 64821 1289
rect 64532 1240 64724 1280
rect 64492 1231 64532 1240
rect 64684 1112 64724 1240
rect 64779 1240 64780 1280
rect 64820 1240 64821 1280
rect 64779 1231 64821 1240
rect 65068 1280 65108 1912
rect 65164 1457 65204 2071
rect 65163 1448 65205 1457
rect 65163 1408 65164 1448
rect 65204 1408 65205 1448
rect 65163 1399 65205 1408
rect 65068 1231 65108 1240
rect 64780 1146 64820 1231
rect 64684 1063 64724 1072
rect 64876 1112 64916 1121
rect 65260 1112 65300 2860
rect 65740 2465 65780 4927
rect 65835 4304 65877 4313
rect 65835 4264 65836 4304
rect 65876 4264 65877 4304
rect 65835 4255 65877 4264
rect 65836 4136 65876 4255
rect 65836 4087 65876 4096
rect 65932 4061 65972 4936
rect 66124 4926 66164 4936
rect 66316 4976 66356 4985
rect 66220 4724 66260 4733
rect 66028 4684 66220 4724
rect 65931 4052 65973 4061
rect 65931 4012 65932 4052
rect 65972 4012 65973 4052
rect 65931 4003 65973 4012
rect 65932 3918 65972 4003
rect 66028 3389 66068 4684
rect 66220 4675 66260 4684
rect 66220 4388 66260 4397
rect 66316 4388 66356 4936
rect 66260 4348 66356 4388
rect 66220 4339 66260 4348
rect 66412 4220 66452 5104
rect 66507 4976 66549 4985
rect 66507 4936 66508 4976
rect 66548 4936 66549 4976
rect 66507 4927 66549 4936
rect 66700 4976 66740 4985
rect 66892 4976 66932 7876
rect 66988 6488 67028 6497
rect 67028 6448 67220 6488
rect 66988 6439 67028 6448
rect 67180 5816 67220 6448
rect 67180 5767 67220 5776
rect 66892 4936 67028 4976
rect 66508 4842 66548 4927
rect 66604 4724 66644 4733
rect 66124 4180 66452 4220
rect 66508 4684 66604 4724
rect 66124 3464 66164 4180
rect 66412 4052 66452 4061
rect 66220 4012 66412 4052
rect 66220 3632 66260 4012
rect 66412 4003 66452 4012
rect 66220 3583 66260 3592
rect 66027 3380 66069 3389
rect 66027 3340 66028 3380
rect 66068 3340 66069 3380
rect 66027 3331 66069 3340
rect 66124 2885 66164 3424
rect 66316 3464 66356 3475
rect 66316 3389 66356 3424
rect 66412 3464 66452 3473
rect 66508 3464 66548 4684
rect 66604 4675 66644 4684
rect 66700 4481 66740 4936
rect 66892 4808 66932 4817
rect 66796 4768 66892 4808
rect 66699 4472 66741 4481
rect 66699 4432 66700 4472
rect 66740 4432 66741 4472
rect 66699 4423 66741 4432
rect 66796 4136 66836 4768
rect 66892 4759 66932 4768
rect 66796 4087 66836 4096
rect 66452 3424 66548 3464
rect 66412 3415 66452 3424
rect 66315 3380 66357 3389
rect 66315 3340 66316 3380
rect 66356 3340 66357 3380
rect 66315 3331 66357 3340
rect 66988 2900 67028 4936
rect 67372 3725 67412 10480
rect 67756 10480 67892 10520
rect 67659 10436 67701 10445
rect 67659 10396 67660 10436
rect 67700 10396 67701 10436
rect 67659 10387 67701 10396
rect 67660 10302 67700 10387
rect 67756 8177 67796 10480
rect 67851 10352 67893 10361
rect 67851 10312 67852 10352
rect 67892 10312 67893 10352
rect 67851 10303 67893 10312
rect 67852 10218 67892 10303
rect 67755 8168 67797 8177
rect 67755 8128 67756 8168
rect 67796 8128 67797 8168
rect 67755 8119 67797 8128
rect 67851 7160 67893 7169
rect 67851 7120 67852 7160
rect 67892 7120 67893 7160
rect 67851 7111 67893 7120
rect 67852 6488 67892 7111
rect 67852 6439 67892 6448
rect 67948 5573 67988 14512
rect 68236 14132 68276 14587
rect 68331 14384 68373 14393
rect 68331 14344 68332 14384
rect 68372 14344 68373 14384
rect 68331 14335 68373 14344
rect 68523 14384 68565 14393
rect 68523 14344 68524 14384
rect 68564 14344 68565 14384
rect 68523 14335 68565 14344
rect 68236 14083 68276 14092
rect 68332 14090 68372 14335
rect 68524 14216 68564 14335
rect 68524 14167 68564 14176
rect 68044 14048 68084 14057
rect 68044 13889 68084 14008
rect 68140 14048 68180 14059
rect 68620 14069 68660 14078
rect 68332 14041 68372 14050
rect 68140 13973 68180 14008
rect 68524 14029 68620 14061
rect 68524 14021 68660 14029
rect 68139 13964 68181 13973
rect 68139 13924 68140 13964
rect 68180 13924 68181 13964
rect 68139 13915 68181 13924
rect 68043 13880 68085 13889
rect 68043 13840 68044 13880
rect 68084 13840 68085 13880
rect 68043 13831 68085 13840
rect 68139 13796 68181 13805
rect 68139 13756 68140 13796
rect 68180 13756 68181 13796
rect 68139 13747 68181 13756
rect 68043 13712 68085 13721
rect 68043 13672 68044 13712
rect 68084 13672 68085 13712
rect 68043 13663 68085 13672
rect 67947 5564 67989 5573
rect 67947 5524 67948 5564
rect 67988 5524 67989 5564
rect 67947 5515 67989 5524
rect 67755 4724 67797 4733
rect 67755 4684 67756 4724
rect 67796 4684 67797 4724
rect 67755 4675 67797 4684
rect 67660 4136 67700 4145
rect 67371 3716 67413 3725
rect 67371 3676 67372 3716
rect 67412 3676 67413 3716
rect 67371 3667 67413 3676
rect 67660 3044 67700 4096
rect 67564 3004 67700 3044
rect 67564 2900 67604 3004
rect 67756 2900 67796 4675
rect 66123 2876 66165 2885
rect 66123 2836 66124 2876
rect 66164 2836 66165 2876
rect 66123 2827 66165 2836
rect 66892 2860 67028 2900
rect 67468 2860 67604 2900
rect 67660 2860 67796 2900
rect 66508 2792 66548 2801
rect 65739 2456 65781 2465
rect 65739 2416 65740 2456
rect 65780 2416 65781 2456
rect 65739 2407 65781 2416
rect 65739 1952 65781 1961
rect 65739 1912 65740 1952
rect 65780 1912 65781 1952
rect 65739 1903 65781 1912
rect 65740 1818 65780 1903
rect 66027 1196 66069 1205
rect 66027 1156 66028 1196
rect 66068 1156 66069 1196
rect 66027 1147 66069 1156
rect 64916 1072 65300 1112
rect 66028 1112 66068 1147
rect 64876 1063 64916 1072
rect 66028 1061 66068 1072
rect 66412 1112 66452 1121
rect 66508 1112 66548 2752
rect 66892 2129 66932 2860
rect 67371 2456 67413 2465
rect 67371 2416 67372 2456
rect 67412 2416 67413 2456
rect 67371 2407 67413 2416
rect 66891 2120 66933 2129
rect 66891 2080 66892 2120
rect 66932 2080 66933 2120
rect 66891 2071 66933 2080
rect 66892 1986 66932 2071
rect 67275 1952 67317 1961
rect 67275 1912 67276 1952
rect 67316 1912 67317 1952
rect 67275 1903 67317 1912
rect 67372 1952 67412 2407
rect 67468 1961 67508 2860
rect 67372 1903 67412 1912
rect 67467 1952 67509 1961
rect 67467 1912 67468 1952
rect 67508 1912 67509 1952
rect 67467 1903 67509 1912
rect 67564 1952 67604 1963
rect 66452 1072 66548 1112
rect 67276 1112 67316 1903
rect 67564 1877 67604 1912
rect 67660 1952 67700 2860
rect 67947 2288 67989 2297
rect 67947 2248 67948 2288
rect 67988 2248 67989 2288
rect 67947 2239 67989 2248
rect 67660 1903 67700 1912
rect 67948 1952 67988 2239
rect 67948 1903 67988 1912
rect 67563 1868 67605 1877
rect 67563 1828 67564 1868
rect 67604 1828 67605 1868
rect 67563 1819 67605 1828
rect 68044 1709 68084 13663
rect 68140 9680 68180 13747
rect 68524 13637 68564 14021
rect 68620 14020 68660 14021
rect 68716 14048 68756 14848
rect 68812 14720 68852 14729
rect 68852 14680 68948 14720
rect 68812 14671 68852 14680
rect 68811 14132 68853 14141
rect 68811 14092 68812 14132
rect 68852 14092 68853 14132
rect 68811 14083 68853 14092
rect 68716 13796 68756 14008
rect 68812 14048 68852 14083
rect 68812 13997 68852 14008
rect 68908 13880 68948 14680
rect 69100 14309 69140 15931
rect 70540 15728 70580 15737
rect 69964 15688 70196 15728
rect 69868 15476 69908 15485
rect 69868 15401 69908 15436
rect 69867 15392 69909 15401
rect 69867 15352 69868 15392
rect 69908 15352 69909 15392
rect 69867 15343 69909 15352
rect 69676 15308 69716 15317
rect 69195 14384 69237 14393
rect 69195 14344 69196 14384
rect 69236 14344 69237 14384
rect 69195 14335 69237 14344
rect 69099 14300 69141 14309
rect 69099 14260 69100 14300
rect 69140 14260 69141 14300
rect 69099 14251 69141 14260
rect 69004 14216 69044 14225
rect 69003 14176 69004 14216
rect 69003 14167 69044 14176
rect 69003 14048 69043 14167
rect 69003 14008 69044 14048
rect 69004 13964 69044 14008
rect 69196 13964 69236 14335
rect 69387 14132 69429 14141
rect 69387 14092 69388 14132
rect 69428 14092 69429 14132
rect 69387 14083 69429 14092
rect 69004 13924 69140 13964
rect 68908 13840 69044 13880
rect 68716 13756 68852 13796
rect 68523 13628 68565 13637
rect 68523 13588 68524 13628
rect 68564 13588 68565 13628
rect 68523 13579 68565 13588
rect 68715 13628 68757 13637
rect 68715 13588 68716 13628
rect 68756 13588 68757 13628
rect 68715 13579 68757 13588
rect 68427 13460 68469 13469
rect 68427 13420 68428 13460
rect 68468 13420 68469 13460
rect 68427 13411 68469 13420
rect 68428 10940 68468 13411
rect 68716 13208 68756 13579
rect 68812 13469 68852 13756
rect 68811 13460 68853 13469
rect 68811 13420 68812 13460
rect 68852 13420 68853 13460
rect 68811 13411 68853 13420
rect 68620 13049 68660 13134
rect 68619 13040 68661 13049
rect 68619 13000 68620 13040
rect 68660 13000 68661 13040
rect 68619 12991 68661 13000
rect 68619 12872 68661 12881
rect 68619 12832 68620 12872
rect 68660 12832 68661 12872
rect 68619 12823 68661 12832
rect 68620 12545 68660 12823
rect 68619 12536 68661 12545
rect 68619 12496 68620 12536
rect 68660 12496 68661 12536
rect 68619 12487 68661 12496
rect 68620 12402 68660 12487
rect 68716 11108 68756 13168
rect 68812 13208 68852 13411
rect 68812 13159 68852 13168
rect 68907 13208 68949 13217
rect 68907 13168 68908 13208
rect 68948 13168 68949 13208
rect 68907 13159 68949 13168
rect 68908 13074 68948 13159
rect 69004 12965 69044 13840
rect 69100 13637 69140 13924
rect 69196 13889 69236 13924
rect 69195 13880 69237 13889
rect 69195 13840 69196 13880
rect 69236 13840 69237 13880
rect 69195 13831 69237 13840
rect 69291 13796 69333 13805
rect 69291 13756 69292 13796
rect 69332 13756 69333 13796
rect 69291 13747 69333 13756
rect 69099 13628 69141 13637
rect 69099 13588 69100 13628
rect 69140 13588 69141 13628
rect 69099 13579 69141 13588
rect 69099 13292 69141 13301
rect 69099 13252 69100 13292
rect 69140 13252 69141 13292
rect 69099 13243 69141 13252
rect 69100 13208 69140 13243
rect 69003 12956 69045 12965
rect 69003 12916 69004 12956
rect 69044 12916 69045 12956
rect 69003 12907 69045 12916
rect 69100 12704 69140 13168
rect 69292 13208 69332 13747
rect 69004 12664 69140 12704
rect 69196 13040 69236 13049
rect 69004 11873 69044 12664
rect 69099 12536 69141 12545
rect 69099 12496 69100 12536
rect 69140 12496 69141 12536
rect 69099 12487 69141 12496
rect 68811 11864 68853 11873
rect 68811 11824 68812 11864
rect 68852 11824 68853 11864
rect 68811 11815 68853 11824
rect 69003 11864 69045 11873
rect 69003 11824 69004 11864
rect 69044 11824 69045 11864
rect 69003 11815 69045 11824
rect 68812 11192 68852 11815
rect 68907 11696 68949 11705
rect 68907 11656 68908 11696
rect 68948 11656 68949 11696
rect 68907 11647 68949 11656
rect 69100 11696 69140 12487
rect 69100 11647 69140 11656
rect 69196 11696 69236 13000
rect 69292 11705 69332 13168
rect 69388 13208 69428 14083
rect 69676 14048 69716 15268
rect 69868 15065 69908 15343
rect 69867 15056 69909 15065
rect 69867 15016 69868 15056
rect 69908 15016 69909 15056
rect 69867 15007 69909 15016
rect 69964 14720 70004 15688
rect 69388 13159 69428 13168
rect 69484 14008 69676 14048
rect 69484 13049 69524 14008
rect 69676 13999 69716 14008
rect 69868 14680 70004 14720
rect 70060 15560 70100 15569
rect 70060 14720 70100 15520
rect 70156 15560 70196 15688
rect 70156 15511 70196 15520
rect 70252 15688 70540 15728
rect 70060 14680 70196 14720
rect 69868 13973 69908 14680
rect 69964 14552 70004 14561
rect 70004 14512 70100 14552
rect 69964 14503 70004 14512
rect 70060 14141 70100 14512
rect 70156 14477 70196 14680
rect 70155 14468 70197 14477
rect 70155 14428 70156 14468
rect 70196 14428 70197 14468
rect 70155 14419 70197 14428
rect 70059 14132 70101 14141
rect 70059 14092 70060 14132
rect 70100 14092 70101 14132
rect 70059 14083 70101 14092
rect 69963 14048 70005 14057
rect 69963 14008 69964 14048
rect 70004 14008 70005 14048
rect 69963 13999 70005 14008
rect 69867 13964 69909 13973
rect 69867 13924 69868 13964
rect 69908 13924 69909 13964
rect 69867 13915 69909 13924
rect 69868 13553 69908 13915
rect 69964 13914 70004 13999
rect 70060 13998 70100 14083
rect 70252 13712 70292 15688
rect 70540 15679 70580 15688
rect 70924 15644 70964 16192
rect 71308 16232 71348 16241
rect 71500 16232 71540 17116
rect 71654 17107 71696 17116
rect 71788 17116 71985 17156
rect 71348 16192 71540 16232
rect 71308 16183 71348 16192
rect 70924 15604 71444 15644
rect 70732 15569 70772 15600
rect 70348 15560 70388 15569
rect 70731 15560 70773 15569
rect 70388 15520 70484 15560
rect 70348 15511 70388 15520
rect 70348 15308 70388 15317
rect 70348 14720 70388 15268
rect 70348 14671 70388 14680
rect 70444 14216 70484 15520
rect 70731 15520 70732 15560
rect 70772 15520 70773 15560
rect 70731 15511 70773 15520
rect 70732 15476 70772 15511
rect 70539 15308 70581 15317
rect 70539 15268 70540 15308
rect 70580 15268 70581 15308
rect 70539 15259 70581 15268
rect 70540 14561 70580 15259
rect 70635 14972 70677 14981
rect 70635 14932 70636 14972
rect 70676 14932 70677 14972
rect 70635 14923 70677 14932
rect 70636 14729 70676 14923
rect 70732 14897 70772 15436
rect 71116 15476 71156 15485
rect 71116 15317 71156 15436
rect 71308 15392 71348 15401
rect 70924 15308 70964 15317
rect 70827 15140 70869 15149
rect 70827 15100 70828 15140
rect 70868 15100 70869 15140
rect 70827 15091 70869 15100
rect 70731 14888 70773 14897
rect 70731 14848 70732 14888
rect 70772 14848 70773 14888
rect 70731 14839 70773 14848
rect 70635 14720 70677 14729
rect 70635 14680 70636 14720
rect 70676 14680 70677 14720
rect 70635 14671 70677 14680
rect 70732 14720 70772 14729
rect 70828 14720 70868 15091
rect 70772 14680 70868 14720
rect 70732 14671 70772 14680
rect 70539 14552 70581 14561
rect 70539 14512 70540 14552
rect 70580 14512 70581 14552
rect 70539 14503 70581 14512
rect 70540 14216 70580 14225
rect 70444 14176 70540 14216
rect 70060 13672 70292 13712
rect 70348 13796 70388 13805
rect 69867 13544 69909 13553
rect 69867 13504 69868 13544
rect 69908 13504 69909 13544
rect 69867 13495 69909 13504
rect 70060 13376 70100 13672
rect 70155 13544 70197 13553
rect 70155 13504 70156 13544
rect 70196 13504 70197 13544
rect 70155 13495 70197 13504
rect 70156 13460 70196 13495
rect 70156 13409 70196 13420
rect 69676 13336 70100 13376
rect 69579 13208 69621 13217
rect 69579 13168 69580 13208
rect 69620 13168 69621 13208
rect 69579 13159 69621 13168
rect 69676 13208 69716 13336
rect 69483 13040 69525 13049
rect 69483 13000 69484 13040
rect 69524 13000 69525 13040
rect 69483 12991 69525 13000
rect 69483 11948 69525 11957
rect 69483 11908 69484 11948
rect 69524 11908 69525 11948
rect 69483 11899 69525 11908
rect 69484 11814 69524 11899
rect 69196 11647 69236 11656
rect 69291 11696 69333 11705
rect 69291 11656 69292 11696
rect 69332 11656 69333 11696
rect 69291 11647 69333 11656
rect 68908 11562 68948 11647
rect 69003 11612 69045 11621
rect 69003 11572 69004 11612
rect 69044 11572 69045 11612
rect 69003 11563 69045 11572
rect 69004 11478 69044 11563
rect 69292 11528 69332 11647
rect 69196 11488 69332 11528
rect 69580 11612 69620 13159
rect 69676 12125 69716 13168
rect 69868 13208 69908 13217
rect 69772 13124 69812 13133
rect 69772 12881 69812 13084
rect 69771 12872 69813 12881
rect 69771 12832 69772 12872
rect 69812 12832 69813 12872
rect 69771 12823 69813 12832
rect 69772 12284 69812 12293
rect 69675 12116 69717 12125
rect 69675 12076 69676 12116
rect 69716 12076 69717 12116
rect 69675 12067 69717 12076
rect 69772 11612 69812 12244
rect 69868 11957 69908 13168
rect 70060 13208 70100 13336
rect 70060 13159 70100 13168
rect 70252 13208 70292 13217
rect 70348 13208 70388 13756
rect 70292 13168 70388 13208
rect 70252 13159 70292 13168
rect 70155 13040 70197 13049
rect 70155 13000 70156 13040
rect 70196 13000 70197 13040
rect 70155 12991 70197 13000
rect 70059 12872 70101 12881
rect 70059 12832 70060 12872
rect 70100 12832 70101 12872
rect 70059 12823 70101 12832
rect 70060 12545 70100 12823
rect 69964 12536 70004 12545
rect 69964 12041 70004 12496
rect 70059 12536 70101 12545
rect 70059 12496 70060 12536
rect 70100 12496 70101 12536
rect 70059 12487 70101 12496
rect 70060 12402 70100 12487
rect 69963 12032 70005 12041
rect 69963 11992 69964 12032
rect 70004 11992 70005 12032
rect 69963 11983 70005 11992
rect 69867 11948 69909 11957
rect 69867 11908 69868 11948
rect 69908 11908 69909 11948
rect 69867 11899 69909 11908
rect 70059 11864 70101 11873
rect 70059 11824 70060 11864
rect 70100 11824 70101 11864
rect 70059 11815 70101 11824
rect 69867 11780 69909 11789
rect 69867 11740 69868 11780
rect 69908 11740 69909 11780
rect 69867 11731 69909 11740
rect 69868 11696 69908 11731
rect 69868 11645 69908 11656
rect 69580 11572 69772 11612
rect 68812 11152 69044 11192
rect 68716 11068 68948 11108
rect 68812 10940 68852 10949
rect 68428 10900 68812 10940
rect 68812 10891 68852 10900
rect 68620 10772 68660 10781
rect 68428 10732 68620 10772
rect 68428 10529 68468 10732
rect 68620 10723 68660 10732
rect 68908 10613 68948 11068
rect 69004 11024 69044 11152
rect 69004 10975 69044 10984
rect 69196 11024 69236 11488
rect 69196 10975 69236 10984
rect 69292 11024 69332 11033
rect 69580 11024 69620 11572
rect 69772 11563 69812 11572
rect 69675 11108 69717 11117
rect 69675 11068 69676 11108
rect 69716 11068 69717 11108
rect 69675 11059 69717 11068
rect 69332 10984 69620 11024
rect 69292 10975 69332 10984
rect 69676 10940 69716 11059
rect 69676 10891 69716 10900
rect 69004 10772 69044 10781
rect 69484 10772 69524 10781
rect 69964 10772 70004 10781
rect 68907 10604 68949 10613
rect 68907 10564 68908 10604
rect 68948 10564 68949 10604
rect 68907 10555 68949 10564
rect 68427 10520 68469 10529
rect 68427 10480 68428 10520
rect 68468 10480 68469 10520
rect 68427 10471 68469 10480
rect 68235 10268 68277 10277
rect 68235 10228 68236 10268
rect 68276 10228 68277 10268
rect 68235 10219 68277 10228
rect 68236 10184 68276 10219
rect 68236 10133 68276 10144
rect 68332 10184 68372 10193
rect 68332 9941 68372 10144
rect 68428 10184 68468 10471
rect 68907 10352 68949 10361
rect 68907 10312 68908 10352
rect 68948 10312 68949 10352
rect 68907 10303 68949 10312
rect 68619 10268 68661 10277
rect 68619 10228 68620 10268
rect 68660 10228 68756 10268
rect 68619 10219 68661 10228
rect 68428 10135 68468 10144
rect 68523 10184 68565 10193
rect 68523 10144 68524 10184
rect 68564 10144 68565 10184
rect 68523 10135 68565 10144
rect 68716 10184 68756 10228
rect 68716 10135 68756 10144
rect 68908 10184 68948 10303
rect 68908 10135 68948 10144
rect 69004 10184 69044 10732
rect 69292 10732 69484 10772
rect 69292 10277 69332 10732
rect 69484 10723 69524 10732
rect 69868 10732 69964 10772
rect 70060 10772 70100 11815
rect 70156 11696 70196 12991
rect 70444 12980 70484 14176
rect 70540 14148 70580 14176
rect 70636 13964 70676 14671
rect 70827 14552 70869 14561
rect 70827 14512 70828 14552
rect 70868 14512 70869 14552
rect 70827 14503 70869 14512
rect 70732 13964 70772 13973
rect 70636 13924 70732 13964
rect 70732 13915 70772 13924
rect 70828 13805 70868 14503
rect 70924 14048 70964 15268
rect 71115 15308 71157 15317
rect 71115 15268 71116 15308
rect 71156 15268 71157 15308
rect 71115 15259 71157 15268
rect 71308 15149 71348 15352
rect 71307 15140 71349 15149
rect 71307 15100 71308 15140
rect 71348 15100 71349 15140
rect 71307 15091 71349 15100
rect 71019 14468 71061 14477
rect 71019 14428 71020 14468
rect 71060 14428 71061 14468
rect 71019 14419 71061 14428
rect 71020 14132 71060 14419
rect 71020 14083 71060 14092
rect 70924 13889 70964 14008
rect 71115 14048 71157 14057
rect 71115 14008 71116 14048
rect 71156 14008 71157 14048
rect 71115 13999 71157 14008
rect 71116 13914 71156 13999
rect 70923 13880 70965 13889
rect 70923 13840 70924 13880
rect 70964 13840 70965 13880
rect 70923 13831 70965 13840
rect 70827 13796 70869 13805
rect 70252 12940 70484 12980
rect 70636 13756 70828 13796
rect 70868 13756 70869 13796
rect 70636 12980 70676 13756
rect 70827 13747 70869 13756
rect 70828 13662 70868 13747
rect 71020 13376 71060 13385
rect 71020 12980 71060 13336
rect 70636 12940 70772 12980
rect 70252 12545 70292 12940
rect 70635 12704 70677 12713
rect 70635 12664 70636 12704
rect 70676 12664 70677 12704
rect 70635 12655 70677 12664
rect 70251 12536 70293 12545
rect 70251 12496 70252 12536
rect 70292 12496 70293 12536
rect 70251 12487 70293 12496
rect 70444 12536 70484 12545
rect 70252 12368 70292 12377
rect 70444 12368 70484 12496
rect 70292 12328 70484 12368
rect 70252 12319 70292 12328
rect 70251 12200 70293 12209
rect 70251 12160 70252 12200
rect 70292 12160 70293 12200
rect 70251 12151 70293 12160
rect 70156 11117 70196 11656
rect 70252 11621 70292 12151
rect 70347 12116 70389 12125
rect 70347 12076 70348 12116
rect 70388 12076 70389 12116
rect 70347 12067 70389 12076
rect 70251 11612 70293 11621
rect 70251 11572 70252 11612
rect 70292 11572 70293 11612
rect 70251 11563 70293 11572
rect 70155 11108 70197 11117
rect 70155 11068 70156 11108
rect 70196 11068 70197 11108
rect 70155 11059 70197 11068
rect 70156 10940 70196 10949
rect 70252 10940 70292 11563
rect 70348 11285 70388 12067
rect 70539 12032 70581 12041
rect 70539 11992 70540 12032
rect 70580 11992 70581 12032
rect 70539 11983 70581 11992
rect 70540 11948 70580 11983
rect 70540 11897 70580 11908
rect 70636 11789 70676 12655
rect 70635 11780 70677 11789
rect 70635 11740 70636 11780
rect 70676 11740 70677 11780
rect 70635 11731 70677 11740
rect 70443 11696 70485 11705
rect 70443 11656 70444 11696
rect 70484 11656 70485 11696
rect 70443 11647 70485 11656
rect 70636 11696 70676 11731
rect 70444 11562 70484 11647
rect 70636 11646 70676 11656
rect 70347 11276 70389 11285
rect 70347 11236 70348 11276
rect 70388 11236 70389 11276
rect 70347 11227 70389 11236
rect 70196 10900 70292 10940
rect 70156 10891 70196 10900
rect 70060 10732 70292 10772
rect 69387 10604 69429 10613
rect 69387 10564 69388 10604
rect 69428 10564 69429 10604
rect 69387 10555 69429 10564
rect 69291 10268 69333 10277
rect 69291 10228 69292 10268
rect 69332 10228 69333 10268
rect 69291 10219 69333 10228
rect 69004 10135 69044 10144
rect 69195 10184 69237 10193
rect 69195 10144 69196 10184
rect 69236 10144 69237 10184
rect 69195 10135 69237 10144
rect 69292 10184 69332 10219
rect 68524 10050 68564 10135
rect 68811 10100 68853 10109
rect 68811 10060 68812 10100
rect 68852 10060 68853 10100
rect 68811 10051 68853 10060
rect 69099 10100 69141 10109
rect 69099 10060 69100 10100
rect 69140 10060 69141 10100
rect 69099 10051 69141 10060
rect 68812 9966 68852 10051
rect 68331 9932 68373 9941
rect 68331 9892 68332 9932
rect 68372 9892 68373 9932
rect 68331 9883 68373 9892
rect 68140 9640 68276 9680
rect 68140 9512 68180 9521
rect 68140 8681 68180 9472
rect 68139 8672 68181 8681
rect 68139 8632 68140 8672
rect 68180 8632 68181 8672
rect 68139 8623 68181 8632
rect 68140 7169 68180 8623
rect 68139 7160 68181 7169
rect 68139 7120 68140 7160
rect 68180 7120 68181 7160
rect 68139 7111 68181 7120
rect 68236 4817 68276 9640
rect 68907 9260 68949 9269
rect 68907 9220 68908 9260
rect 68948 9220 68949 9260
rect 68907 9211 68949 9220
rect 68524 8840 68564 8849
rect 68427 8336 68469 8345
rect 68427 8296 68428 8336
rect 68468 8296 68469 8336
rect 68427 8287 68469 8296
rect 68428 8168 68468 8287
rect 68428 8119 68468 8128
rect 68524 7916 68564 8800
rect 68715 8672 68757 8681
rect 68715 8632 68716 8672
rect 68756 8632 68757 8672
rect 68715 8623 68757 8632
rect 68908 8672 68948 9211
rect 69003 8840 69045 8849
rect 69003 8800 69004 8840
rect 69044 8800 69045 8840
rect 69003 8791 69045 8800
rect 68908 8623 68948 8632
rect 69004 8672 69044 8791
rect 69004 8623 69044 8632
rect 68716 8538 68756 8623
rect 68812 8504 68852 8513
rect 68620 8084 68660 8093
rect 68812 8084 68852 8464
rect 68660 8044 68852 8084
rect 68620 8035 68660 8044
rect 69004 8000 69044 8009
rect 68716 7960 69004 8000
rect 68716 7916 68756 7960
rect 69004 7951 69044 7960
rect 68524 7876 68756 7916
rect 68427 7748 68469 7757
rect 68427 7708 68428 7748
rect 68468 7708 68469 7748
rect 68427 7699 68469 7708
rect 68428 7614 68468 7699
rect 69100 7085 69140 10051
rect 69196 9680 69236 10135
rect 69292 10134 69332 10144
rect 69292 9680 69332 9689
rect 69196 9640 69292 9680
rect 69292 9631 69332 9640
rect 69388 9437 69428 10555
rect 69483 10520 69525 10529
rect 69483 10480 69484 10520
rect 69524 10480 69525 10520
rect 69483 10471 69525 10480
rect 69484 9596 69524 10471
rect 69771 10352 69813 10361
rect 69771 10312 69772 10352
rect 69812 10312 69813 10352
rect 69771 10303 69813 10312
rect 69580 10184 69620 10195
rect 69580 10109 69620 10144
rect 69675 10184 69717 10193
rect 69675 10144 69676 10184
rect 69716 10144 69717 10184
rect 69675 10135 69717 10144
rect 69579 10100 69621 10109
rect 69579 10060 69580 10100
rect 69620 10060 69621 10100
rect 69579 10051 69621 10060
rect 69676 10050 69716 10135
rect 69675 9932 69717 9941
rect 69675 9892 69676 9932
rect 69716 9892 69717 9932
rect 69675 9883 69717 9892
rect 69676 9680 69716 9883
rect 69676 9631 69716 9640
rect 69484 9556 69620 9596
rect 69387 9428 69429 9437
rect 69474 9428 69514 9434
rect 69387 9388 69388 9428
rect 69428 9425 69514 9428
rect 69428 9388 69474 9425
rect 69387 9379 69429 9388
rect 69474 9376 69514 9385
rect 69292 9260 69332 9269
rect 69332 9220 69524 9260
rect 69292 9211 69332 9220
rect 69291 9008 69333 9017
rect 69291 8968 69292 9008
rect 69332 8968 69333 9008
rect 69291 8959 69333 8968
rect 69196 8849 69236 8934
rect 69195 8840 69237 8849
rect 69195 8800 69196 8840
rect 69236 8800 69237 8840
rect 69195 8791 69237 8800
rect 69196 8672 69236 8683
rect 69196 8597 69236 8632
rect 69195 8588 69237 8597
rect 69195 8548 69196 8588
rect 69236 8548 69237 8588
rect 69195 8539 69237 8548
rect 69292 7496 69332 8959
rect 69387 8840 69429 8849
rect 69387 8800 69388 8840
rect 69428 8800 69429 8840
rect 69387 8791 69429 8800
rect 69388 8672 69428 8791
rect 69388 8623 69428 8632
rect 69484 8672 69524 9220
rect 69580 8840 69620 9556
rect 69676 9260 69716 9269
rect 69676 9017 69716 9220
rect 69675 9008 69717 9017
rect 69675 8968 69676 9008
rect 69716 8968 69717 9008
rect 69675 8959 69717 8968
rect 69772 8924 69812 10303
rect 69868 9605 69908 10732
rect 69964 10723 70004 10732
rect 69964 10352 70004 10361
rect 69867 9596 69909 9605
rect 69867 9556 69868 9596
rect 69908 9556 69909 9596
rect 69867 9547 69909 9556
rect 69868 9512 69908 9547
rect 69868 9462 69908 9472
rect 69867 9344 69909 9353
rect 69867 9304 69868 9344
rect 69908 9304 69909 9344
rect 69867 9295 69909 9304
rect 69868 9210 69908 9295
rect 69772 8875 69812 8884
rect 69580 8800 69716 8840
rect 69676 8756 69716 8800
rect 69676 8716 69812 8756
rect 69484 8623 69524 8632
rect 69579 8672 69621 8681
rect 69579 8632 69580 8672
rect 69620 8632 69621 8672
rect 69579 8623 69621 8632
rect 69676 8651 69716 8660
rect 69292 7456 69524 7496
rect 69388 7328 69428 7337
rect 69099 7076 69141 7085
rect 69099 7036 69100 7076
rect 69140 7036 69141 7076
rect 69099 7027 69141 7036
rect 69004 6656 69044 6665
rect 69100 6656 69140 7027
rect 69044 6616 69140 6656
rect 69004 6607 69044 6616
rect 69196 6488 69236 6497
rect 69388 6488 69428 7288
rect 69484 6992 69524 7456
rect 69580 7160 69620 8623
rect 69676 8513 69716 8611
rect 69675 8504 69717 8513
rect 69675 8464 69676 8504
rect 69716 8464 69717 8504
rect 69675 8455 69717 8464
rect 69580 7111 69620 7120
rect 69676 7160 69716 7169
rect 69676 6992 69716 7120
rect 69484 6952 69716 6992
rect 69580 6488 69620 6497
rect 69388 6448 69580 6488
rect 69196 5909 69236 6448
rect 69580 6439 69620 6448
rect 69387 6068 69429 6077
rect 69387 6028 69388 6068
rect 69428 6028 69429 6068
rect 69387 6019 69429 6028
rect 69195 5900 69237 5909
rect 69195 5860 69196 5900
rect 69236 5860 69237 5900
rect 69195 5851 69237 5860
rect 69099 5648 69141 5657
rect 69099 5608 69100 5648
rect 69140 5608 69141 5648
rect 69099 5599 69141 5608
rect 69291 5648 69333 5657
rect 69291 5599 69292 5648
rect 68812 4976 68852 4985
rect 69004 4976 69044 4985
rect 68852 4936 68948 4976
rect 68812 4927 68852 4936
rect 68235 4808 68277 4817
rect 68235 4768 68236 4808
rect 68276 4768 68277 4808
rect 68235 4759 68277 4768
rect 68811 4724 68853 4733
rect 68811 4684 68812 4724
rect 68852 4684 68853 4724
rect 68811 4675 68853 4684
rect 68812 4590 68852 4675
rect 68811 4472 68853 4481
rect 68811 4432 68812 4472
rect 68852 4432 68853 4472
rect 68811 4423 68853 4432
rect 68715 4304 68757 4313
rect 68715 4264 68716 4304
rect 68756 4264 68757 4304
rect 68715 4255 68757 4264
rect 68812 4304 68852 4423
rect 68812 4255 68852 4264
rect 68620 3464 68660 3473
rect 68235 3296 68277 3305
rect 68235 3256 68236 3296
rect 68276 3256 68277 3296
rect 68235 3247 68277 3256
rect 68236 2624 68276 3247
rect 68620 2900 68660 3424
rect 68716 3464 68756 4255
rect 68811 4136 68853 4145
rect 68811 4096 68812 4136
rect 68852 4096 68853 4136
rect 68811 4087 68853 4096
rect 68716 3137 68756 3424
rect 68715 3128 68757 3137
rect 68715 3088 68716 3128
rect 68756 3088 68757 3128
rect 68715 3079 68757 3088
rect 68428 2860 68660 2900
rect 68236 2575 68276 2584
rect 68332 2624 68372 2635
rect 68332 2549 68372 2584
rect 68428 2624 68468 2860
rect 68716 2792 68756 2801
rect 68331 2540 68373 2549
rect 68331 2500 68332 2540
rect 68372 2500 68373 2540
rect 68331 2491 68373 2500
rect 68139 2456 68181 2465
rect 68139 2416 68140 2456
rect 68180 2416 68181 2456
rect 68139 2407 68181 2416
rect 68140 2322 68180 2407
rect 68235 2372 68277 2381
rect 68235 2332 68236 2372
rect 68276 2332 68277 2372
rect 68235 2323 68277 2332
rect 68236 1952 68276 2323
rect 68236 1903 68276 1912
rect 68332 1952 68372 1961
rect 68428 1952 68468 2584
rect 68372 1912 68468 1952
rect 68332 1903 68372 1912
rect 67372 1700 67412 1709
rect 67372 1205 67412 1660
rect 68043 1700 68085 1709
rect 68043 1660 68044 1700
rect 68084 1660 68085 1700
rect 68043 1651 68085 1660
rect 68428 1364 68468 1912
rect 68524 2752 68716 2792
rect 68524 1877 68564 2752
rect 68716 2743 68756 2752
rect 68620 2624 68660 2633
rect 68523 1868 68565 1877
rect 68523 1828 68524 1868
rect 68564 1828 68565 1868
rect 68523 1819 68565 1828
rect 68428 1315 68468 1324
rect 67371 1196 67413 1205
rect 67371 1156 67372 1196
rect 67412 1156 67413 1196
rect 67371 1147 67413 1156
rect 66412 1063 66452 1072
rect 67276 1063 67316 1072
rect 64204 953 64244 988
rect 58923 944 58965 953
rect 58923 904 58924 944
rect 58964 904 58965 944
rect 58923 895 58965 904
rect 60363 944 60405 953
rect 60363 904 60364 944
rect 60404 904 60405 944
rect 60363 895 60405 904
rect 62955 944 62997 953
rect 62955 904 62956 944
rect 62996 904 62997 944
rect 62955 895 62997 904
rect 63723 944 63765 953
rect 63723 904 63724 944
rect 63764 904 63765 944
rect 63723 895 63765 904
rect 64203 944 64245 953
rect 64203 904 64204 944
rect 64244 904 64245 944
rect 68524 944 68564 1819
rect 68620 1784 68660 2584
rect 68812 2624 68852 4087
rect 68908 3473 68948 4936
rect 69004 4313 69044 4936
rect 69100 4976 69140 5599
rect 69332 5599 69333 5648
rect 69388 5648 69428 6019
rect 69676 5816 69716 6952
rect 69772 7160 69812 8716
rect 69868 8672 69908 8681
rect 69964 8672 70004 10312
rect 70059 10352 70101 10361
rect 70059 10312 70060 10352
rect 70100 10312 70101 10352
rect 70059 10303 70101 10312
rect 70060 9512 70100 10303
rect 70060 9463 70100 9472
rect 70155 9512 70197 9521
rect 70155 9472 70156 9512
rect 70196 9472 70197 9512
rect 70155 9463 70197 9472
rect 70156 9378 70196 9463
rect 69908 8632 70004 8672
rect 70060 8840 70100 8849
rect 69868 8623 69908 8632
rect 70060 8597 70100 8800
rect 70155 8840 70197 8849
rect 70155 8800 70156 8840
rect 70196 8800 70197 8840
rect 70155 8791 70197 8800
rect 70059 8588 70101 8597
rect 70059 8548 70060 8588
rect 70100 8548 70101 8588
rect 70059 8539 70101 8548
rect 69868 8000 69908 8009
rect 69908 7960 70004 8000
rect 69868 7951 69908 7960
rect 69867 7244 69909 7253
rect 69867 7204 69868 7244
rect 69908 7204 69909 7244
rect 69867 7195 69909 7204
rect 69772 6077 69812 7120
rect 69868 7160 69908 7195
rect 69964 7169 70004 7960
rect 69868 7109 69908 7120
rect 69963 7160 70005 7169
rect 69963 7120 69964 7160
rect 70004 7120 70005 7160
rect 69963 7111 70005 7120
rect 70060 7160 70100 8539
rect 70156 7328 70196 8791
rect 70252 8756 70292 10732
rect 70348 9428 70388 11227
rect 70540 10940 70580 10949
rect 70732 10940 70772 12940
rect 70828 12940 71060 12980
rect 70828 12536 70868 12940
rect 70828 12487 70868 12496
rect 70580 10900 70772 10940
rect 71116 10940 71156 10949
rect 70540 10891 70580 10900
rect 71116 10781 71156 10900
rect 71308 10856 71348 10865
rect 70731 10772 70773 10781
rect 70731 10732 70732 10772
rect 70772 10732 70773 10772
rect 70731 10723 70773 10732
rect 70924 10772 70964 10781
rect 70732 10638 70772 10723
rect 70924 10352 70964 10732
rect 71115 10772 71157 10781
rect 71115 10732 71116 10772
rect 71156 10732 71157 10772
rect 71115 10723 71157 10732
rect 70732 10312 70964 10352
rect 70635 10268 70677 10277
rect 70635 10228 70636 10268
rect 70676 10228 70677 10268
rect 70635 10219 70677 10228
rect 70348 9379 70388 9388
rect 70444 10100 70484 10109
rect 70444 9353 70484 10060
rect 70443 9344 70485 9353
rect 70443 9304 70444 9344
rect 70484 9304 70485 9344
rect 70443 9295 70485 9304
rect 70540 9260 70580 9269
rect 70540 9101 70580 9220
rect 70539 9092 70581 9101
rect 70252 8707 70292 8716
rect 70444 9052 70540 9092
rect 70580 9052 70581 9092
rect 70444 8651 70484 9052
rect 70539 9043 70581 9052
rect 70636 8672 70676 10219
rect 70732 9512 70772 10312
rect 70827 10184 70869 10193
rect 70827 10144 70828 10184
rect 70868 10144 70869 10184
rect 70827 10135 70869 10144
rect 70828 10050 70868 10135
rect 70923 10016 70965 10025
rect 70923 9976 70924 10016
rect 70964 9976 70965 10016
rect 70923 9967 70965 9976
rect 70732 8849 70772 9472
rect 70827 9512 70869 9521
rect 70827 9472 70828 9512
rect 70868 9472 70869 9512
rect 70827 9463 70869 9472
rect 70924 9512 70964 9967
rect 71116 9941 71156 10723
rect 71308 10193 71348 10816
rect 71307 10184 71349 10193
rect 71307 10144 71308 10184
rect 71348 10144 71349 10184
rect 71307 10135 71349 10144
rect 71115 9932 71157 9941
rect 71115 9892 71116 9932
rect 71156 9892 71157 9932
rect 71115 9883 71157 9892
rect 71404 9764 71444 15604
rect 71500 10445 71540 16192
rect 71788 16232 71828 17116
rect 72055 17072 72095 17472
rect 72345 17156 72385 17472
rect 71884 17032 72095 17072
rect 72172 17116 72385 17156
rect 71884 16484 71924 17032
rect 71884 16435 71924 16444
rect 71596 14720 71636 14729
rect 71596 12965 71636 14680
rect 71595 12956 71637 12965
rect 71595 12916 71596 12956
rect 71636 12916 71637 12956
rect 71595 12907 71637 12916
rect 71596 12536 71636 12907
rect 71788 12797 71828 16192
rect 72172 16232 72212 17116
rect 72455 17072 72495 17472
rect 72745 17156 72785 17472
rect 72268 17032 72495 17072
rect 72556 17116 72785 17156
rect 72268 16484 72308 17032
rect 72268 16435 72308 16444
rect 71979 16148 72021 16157
rect 71979 16108 71980 16148
rect 72020 16108 72021 16148
rect 71979 16099 72021 16108
rect 71980 13544 72020 16099
rect 72172 15233 72212 16192
rect 72556 16232 72596 17116
rect 72855 17072 72895 17472
rect 73145 17156 73185 17472
rect 72652 17032 72895 17072
rect 72940 17116 73185 17156
rect 72652 16484 72692 17032
rect 72652 16435 72692 16444
rect 72940 16232 72980 17116
rect 73255 17072 73295 17472
rect 73545 17240 73585 17472
rect 73036 17032 73295 17072
rect 73420 17200 73585 17240
rect 73036 16484 73076 17032
rect 73420 16988 73460 17200
rect 73655 17072 73695 17472
rect 73945 17156 73985 17472
rect 73036 16435 73076 16444
rect 73324 16948 73460 16988
rect 73516 17032 73695 17072
rect 73900 17116 73985 17156
rect 72556 15737 72596 16192
rect 72748 16192 72940 16232
rect 72555 15728 72597 15737
rect 72555 15688 72556 15728
rect 72596 15688 72597 15728
rect 72555 15679 72597 15688
rect 72652 15392 72692 15401
rect 72171 15224 72213 15233
rect 72171 15184 72172 15224
rect 72212 15184 72213 15224
rect 72171 15175 72213 15184
rect 72171 14552 72213 14561
rect 72171 14512 72172 14552
rect 72212 14512 72213 14552
rect 72171 14503 72213 14512
rect 72172 14132 72212 14503
rect 72172 14083 72212 14092
rect 72556 14048 72596 14057
rect 72652 14048 72692 15352
rect 72748 14972 72788 16192
rect 72940 16183 72980 16192
rect 73324 16232 73364 16948
rect 73420 16484 73460 16493
rect 73516 16484 73556 17032
rect 73460 16444 73556 16484
rect 73420 16416 73460 16444
rect 73708 16232 73748 16241
rect 73900 16232 73940 17116
rect 74055 17072 74095 17472
rect 74345 17156 74385 17472
rect 72748 14923 72788 14932
rect 72748 14552 72788 14561
rect 72748 14057 72788 14512
rect 72596 14008 72692 14048
rect 72747 14048 72789 14057
rect 72747 14008 72748 14048
rect 72788 14008 72789 14048
rect 72556 13999 72596 14008
rect 72747 13999 72789 14008
rect 71884 13504 72020 13544
rect 71884 13208 71924 13504
rect 71980 13376 72020 13385
rect 72020 13336 72308 13376
rect 71980 13327 72020 13336
rect 72171 13208 72213 13217
rect 71884 13168 72020 13208
rect 71787 12788 71829 12797
rect 71787 12748 71788 12788
rect 71828 12748 71829 12788
rect 71787 12739 71829 12748
rect 71692 12536 71732 12545
rect 71596 12496 71692 12536
rect 71692 12487 71732 12496
rect 71499 10436 71541 10445
rect 71499 10396 71500 10436
rect 71540 10396 71541 10436
rect 71499 10387 71541 10396
rect 71691 10184 71733 10193
rect 71691 10144 71692 10184
rect 71732 10144 71733 10184
rect 71691 10135 71733 10144
rect 71692 10050 71732 10135
rect 71691 9932 71733 9941
rect 71691 9892 71692 9932
rect 71732 9892 71733 9932
rect 71691 9883 71733 9892
rect 70924 9463 70964 9472
rect 71020 9724 71444 9764
rect 70828 9378 70868 9463
rect 70731 8840 70773 8849
rect 70731 8800 70732 8840
rect 70772 8800 70773 8840
rect 70731 8791 70773 8800
rect 70828 8672 70868 8681
rect 70348 8611 70517 8651
rect 70636 8632 70828 8672
rect 70348 8513 70388 8611
rect 70477 8588 70517 8611
rect 70477 8548 70676 8588
rect 70347 8504 70389 8513
rect 70347 8464 70348 8504
rect 70388 8464 70389 8504
rect 70347 8455 70389 8464
rect 70347 7748 70389 7757
rect 70347 7708 70348 7748
rect 70388 7708 70389 7748
rect 70347 7699 70389 7708
rect 70156 7288 70292 7328
rect 70155 7160 70197 7169
rect 70100 7120 70156 7160
rect 70196 7120 70197 7160
rect 70060 7111 70100 7120
rect 70155 7111 70197 7120
rect 70252 7160 70292 7288
rect 70348 7253 70388 7699
rect 70347 7244 70389 7253
rect 70347 7204 70348 7244
rect 70388 7204 70389 7244
rect 70347 7195 70389 7204
rect 69964 6497 70004 7111
rect 70156 6992 70196 7001
rect 70060 6952 70156 6992
rect 69963 6488 70005 6497
rect 69963 6448 69964 6488
rect 70004 6448 70005 6488
rect 69963 6439 70005 6448
rect 69771 6068 69813 6077
rect 69771 6028 69772 6068
rect 69812 6028 69908 6068
rect 69771 6019 69813 6028
rect 69771 5900 69813 5909
rect 69771 5860 69772 5900
rect 69812 5860 69813 5900
rect 69771 5851 69813 5860
rect 69388 5599 69428 5608
rect 69484 5776 69716 5816
rect 69484 5648 69524 5776
rect 69772 5766 69812 5851
rect 69292 5513 69332 5587
rect 69484 5480 69524 5608
rect 69580 5648 69620 5657
rect 69772 5648 69812 5657
rect 69620 5608 69772 5648
rect 69580 5599 69620 5608
rect 69772 5599 69812 5608
rect 69484 5440 69812 5480
rect 69100 4927 69140 4936
rect 69484 4808 69524 4817
rect 69388 4768 69484 4808
rect 69195 4724 69237 4733
rect 69195 4684 69196 4724
rect 69236 4684 69237 4724
rect 69195 4675 69237 4684
rect 69003 4304 69045 4313
rect 69003 4264 69004 4304
rect 69044 4264 69045 4304
rect 69003 4255 69045 4264
rect 69004 4052 69044 4061
rect 69004 3641 69044 4012
rect 69003 3632 69045 3641
rect 69003 3592 69004 3632
rect 69044 3592 69045 3632
rect 69003 3583 69045 3592
rect 68907 3464 68949 3473
rect 68907 3424 68908 3464
rect 68948 3424 68949 3464
rect 68907 3415 68949 3424
rect 69100 3464 69140 3473
rect 68908 3296 68948 3305
rect 69100 3296 69140 3424
rect 69196 3464 69236 4675
rect 69388 4136 69428 4768
rect 69484 4759 69524 4768
rect 69388 4087 69428 4096
rect 69291 3632 69333 3641
rect 69291 3592 69292 3632
rect 69332 3592 69333 3632
rect 69291 3583 69333 3592
rect 69292 3498 69332 3583
rect 69196 3415 69236 3424
rect 69388 3464 69428 3473
rect 69676 3464 69716 3473
rect 69428 3424 69676 3464
rect 69388 3415 69428 3424
rect 69676 3415 69716 3424
rect 69772 3464 69812 5440
rect 69772 3305 69812 3424
rect 69868 3464 69908 6028
rect 69963 5648 70005 5657
rect 69963 5608 69964 5648
rect 70004 5608 70005 5648
rect 69963 5599 70005 5608
rect 70060 5648 70100 6952
rect 70156 6943 70196 6952
rect 70060 5599 70100 5608
rect 69964 5514 70004 5599
rect 70252 4313 70292 7120
rect 70348 7160 70388 7195
rect 70348 7110 70388 7120
rect 70539 7160 70581 7169
rect 70539 7120 70540 7160
rect 70580 7120 70581 7160
rect 70539 7111 70581 7120
rect 70443 6488 70485 6497
rect 70443 6448 70444 6488
rect 70484 6448 70485 6488
rect 70443 6439 70485 6448
rect 70444 6354 70484 6439
rect 70443 4388 70485 4397
rect 70443 4348 70444 4388
rect 70484 4348 70485 4388
rect 70443 4339 70485 4348
rect 70251 4304 70293 4313
rect 70251 4264 70252 4304
rect 70292 4264 70293 4304
rect 70251 4255 70293 4264
rect 70444 4145 70484 4339
rect 70252 4136 70292 4145
rect 69963 3548 70005 3557
rect 69963 3508 69964 3548
rect 70004 3508 70005 3548
rect 69963 3499 70005 3508
rect 68948 3256 69140 3296
rect 69771 3296 69813 3305
rect 69771 3256 69772 3296
rect 69812 3256 69813 3296
rect 68908 3247 68948 3256
rect 69771 3247 69813 3256
rect 69003 3128 69045 3137
rect 69003 3088 69004 3128
rect 69044 3088 69045 3128
rect 69003 3079 69045 3088
rect 68812 2575 68852 2584
rect 69004 2624 69044 3079
rect 69004 2575 69044 2584
rect 69196 2624 69236 2633
rect 69100 2540 69140 2549
rect 69100 2120 69140 2500
rect 69196 2381 69236 2584
rect 69868 2549 69908 3424
rect 69964 3464 70004 3499
rect 70252 3473 70292 4096
rect 70443 4136 70485 4145
rect 70443 4096 70444 4136
rect 70484 4096 70485 4136
rect 70443 4087 70485 4096
rect 69964 3413 70004 3424
rect 70251 3464 70293 3473
rect 70251 3424 70252 3464
rect 70292 3424 70293 3464
rect 70251 3415 70293 3424
rect 69867 2540 69909 2549
rect 69867 2500 69868 2540
rect 69908 2500 69909 2540
rect 69867 2491 69909 2500
rect 69195 2372 69237 2381
rect 69195 2332 69196 2372
rect 69236 2332 69237 2372
rect 69195 2323 69237 2332
rect 68620 1735 68660 1744
rect 68716 2080 69140 2120
rect 68716 1616 68756 2080
rect 70252 1961 70292 3415
rect 70540 3389 70580 7111
rect 70636 4397 70676 8548
rect 70828 5657 70868 8632
rect 71020 8345 71060 9724
rect 71211 9596 71253 9605
rect 71211 9556 71212 9596
rect 71252 9556 71253 9596
rect 71211 9547 71253 9556
rect 71115 9512 71157 9521
rect 71115 9472 71116 9512
rect 71156 9472 71157 9512
rect 71115 9463 71157 9472
rect 71116 8672 71156 9463
rect 71212 8756 71252 9547
rect 71308 9512 71348 9521
rect 71308 9185 71348 9472
rect 71500 9512 71540 9521
rect 71403 9260 71445 9269
rect 71403 9220 71404 9260
rect 71444 9220 71445 9260
rect 71403 9211 71445 9220
rect 71307 9176 71349 9185
rect 71307 9136 71308 9176
rect 71348 9136 71349 9176
rect 71307 9127 71349 9136
rect 71404 9126 71444 9211
rect 71500 8924 71540 9472
rect 71692 9512 71732 9883
rect 71692 9437 71732 9472
rect 71883 9512 71925 9521
rect 71883 9472 71884 9512
rect 71924 9472 71925 9512
rect 71883 9463 71925 9472
rect 71691 9428 71733 9437
rect 71691 9388 71692 9428
rect 71732 9388 71733 9428
rect 71691 9379 71733 9388
rect 71884 9378 71924 9463
rect 71500 8875 71540 8884
rect 71788 9260 71828 9269
rect 71212 8716 71444 8756
rect 71116 8623 71156 8632
rect 71212 8588 71252 8597
rect 71019 8336 71061 8345
rect 71019 8296 71020 8336
rect 71060 8296 71061 8336
rect 71019 8287 71061 8296
rect 71020 8168 71060 8177
rect 71212 8168 71252 8548
rect 71060 8128 71252 8168
rect 71020 8119 71060 8128
rect 71404 8000 71444 8716
rect 71692 8588 71732 8597
rect 71500 8548 71692 8588
rect 71500 8168 71540 8548
rect 71692 8539 71732 8548
rect 71500 8119 71540 8128
rect 71019 7748 71061 7757
rect 71019 7708 71020 7748
rect 71060 7708 71061 7748
rect 71019 7699 71061 7708
rect 71020 7614 71060 7699
rect 71404 7160 71444 7960
rect 71596 8000 71636 8009
rect 71596 7832 71636 7960
rect 71692 8000 71732 8009
rect 71788 8000 71828 9220
rect 71883 9260 71925 9269
rect 71883 9220 71884 9260
rect 71924 9220 71925 9260
rect 71883 9211 71925 9220
rect 71732 7960 71828 8000
rect 71692 7951 71732 7960
rect 71884 7832 71924 9211
rect 71596 7792 71924 7832
rect 71980 7664 72020 13168
rect 72171 13168 72172 13208
rect 72212 13168 72213 13208
rect 72268 13208 72308 13336
rect 72556 13208 72596 13217
rect 72268 13168 72556 13208
rect 72171 13159 72213 13168
rect 72556 13159 72596 13168
rect 72172 13074 72212 13159
rect 73035 12956 73077 12965
rect 73035 12916 73036 12956
rect 73076 12916 73077 12956
rect 73035 12907 73077 12916
rect 72843 12704 72885 12713
rect 72843 12664 72844 12704
rect 72884 12664 72885 12704
rect 72843 12655 72885 12664
rect 72844 12570 72884 12655
rect 72844 11696 72884 11705
rect 72884 11656 72980 11696
rect 72844 11647 72884 11656
rect 72460 11612 72500 11621
rect 72460 11201 72500 11572
rect 72459 11192 72501 11201
rect 72459 11152 72460 11192
rect 72500 11152 72501 11192
rect 72459 11143 72501 11152
rect 72940 10856 72980 11656
rect 72940 10807 72980 10816
rect 72843 10436 72885 10445
rect 72843 10396 72844 10436
rect 72884 10396 72885 10436
rect 72843 10387 72885 10396
rect 72844 10109 72884 10387
rect 72939 10184 72981 10193
rect 72939 10144 72940 10184
rect 72980 10144 72981 10184
rect 72939 10135 72981 10144
rect 72843 10100 72885 10109
rect 72843 10060 72844 10100
rect 72884 10060 72885 10100
rect 72843 10051 72885 10060
rect 72555 9764 72597 9773
rect 72555 9724 72556 9764
rect 72596 9724 72597 9764
rect 72555 9715 72597 9724
rect 72556 9437 72596 9715
rect 72555 9428 72597 9437
rect 72555 9388 72556 9428
rect 72596 9388 72597 9428
rect 72555 9379 72597 9388
rect 72172 9344 72212 9353
rect 72076 9304 72172 9344
rect 72076 8672 72116 9304
rect 72172 9295 72212 9304
rect 72076 8623 72116 8632
rect 71980 7624 72116 7664
rect 71692 7160 71732 7169
rect 71404 7120 71692 7160
rect 70827 5648 70869 5657
rect 70827 5608 70828 5648
rect 70868 5608 70869 5648
rect 70827 5599 70869 5608
rect 71307 5648 71349 5657
rect 71307 5608 71308 5648
rect 71348 5608 71349 5648
rect 71307 5599 71349 5608
rect 71308 5514 71348 5599
rect 71500 4985 71540 7120
rect 71692 7111 71732 7120
rect 71884 7160 71924 7169
rect 71788 6992 71828 7001
rect 71788 6833 71828 6952
rect 71787 6824 71829 6833
rect 71787 6784 71788 6824
rect 71828 6784 71829 6824
rect 71787 6775 71829 6784
rect 71884 6656 71924 7120
rect 71979 7160 72021 7169
rect 71979 7120 71980 7160
rect 72020 7120 72021 7160
rect 71979 7111 72021 7120
rect 71980 7026 72020 7111
rect 71979 6824 72021 6833
rect 71979 6784 71980 6824
rect 72020 6784 72021 6824
rect 71979 6775 72021 6784
rect 71788 6616 71924 6656
rect 71596 6236 71636 6245
rect 71636 6196 71732 6236
rect 71596 6187 71636 6196
rect 71692 5741 71732 6196
rect 71691 5732 71733 5741
rect 71691 5692 71692 5732
rect 71732 5692 71733 5732
rect 71691 5683 71733 5692
rect 71595 5648 71637 5657
rect 71595 5608 71596 5648
rect 71636 5608 71637 5648
rect 71595 5599 71637 5608
rect 71692 5648 71732 5683
rect 71596 5514 71636 5599
rect 71692 5598 71732 5608
rect 71788 5573 71828 6616
rect 71980 6572 72020 6775
rect 71980 6523 72020 6532
rect 71883 6488 71925 6497
rect 71883 6448 71884 6488
rect 71924 6448 71925 6488
rect 71883 6439 71925 6448
rect 71884 5648 71924 6439
rect 71980 5825 72020 5910
rect 71979 5816 72021 5825
rect 71979 5776 71980 5816
rect 72020 5776 72021 5816
rect 71979 5767 72021 5776
rect 71884 5608 72020 5648
rect 71787 5564 71829 5573
rect 71787 5524 71788 5564
rect 71828 5524 71829 5564
rect 71787 5515 71829 5524
rect 70827 4976 70869 4985
rect 71212 4976 71252 4985
rect 70827 4936 70828 4976
rect 70868 4936 70869 4976
rect 70827 4927 70869 4936
rect 71116 4936 71212 4976
rect 70635 4388 70677 4397
rect 70635 4348 70636 4388
rect 70676 4348 70677 4388
rect 70635 4339 70677 4348
rect 70731 4304 70773 4313
rect 70731 4264 70732 4304
rect 70772 4264 70773 4304
rect 70731 4255 70773 4264
rect 70732 3641 70772 4255
rect 70731 3632 70773 3641
rect 70731 3592 70732 3632
rect 70772 3592 70773 3632
rect 70731 3583 70773 3592
rect 70635 3548 70677 3557
rect 70635 3508 70636 3548
rect 70676 3508 70677 3548
rect 70635 3499 70677 3508
rect 70636 3464 70676 3499
rect 70636 3413 70676 3424
rect 70732 3464 70772 3583
rect 70732 3415 70772 3424
rect 70539 3380 70581 3389
rect 70539 3340 70540 3380
rect 70580 3340 70581 3380
rect 70539 3331 70581 3340
rect 68620 1576 68756 1616
rect 68812 1952 68852 1961
rect 68620 1112 68660 1576
rect 68812 1364 68852 1912
rect 69196 1952 69236 1961
rect 70059 1952 70101 1961
rect 69236 1912 69428 1952
rect 69196 1903 69236 1912
rect 69003 1868 69045 1877
rect 69003 1828 69004 1868
rect 69044 1828 69045 1868
rect 69003 1819 69045 1828
rect 68908 1364 68948 1373
rect 68812 1324 68908 1364
rect 68908 1315 68948 1324
rect 68620 1063 68660 1072
rect 68716 1112 68756 1121
rect 68716 944 68756 1072
rect 68908 1112 68948 1121
rect 69004 1112 69044 1819
rect 69388 1280 69428 1912
rect 70059 1912 70060 1952
rect 70100 1912 70101 1952
rect 70059 1903 70101 1912
rect 70251 1952 70293 1961
rect 70251 1912 70252 1952
rect 70292 1912 70293 1952
rect 70251 1903 70293 1912
rect 70060 1364 70100 1903
rect 70828 1877 70868 4927
rect 70924 3464 70964 3475
rect 70924 3389 70964 3424
rect 70923 3380 70965 3389
rect 70923 3340 70924 3380
rect 70964 3340 70965 3380
rect 70923 3331 70965 3340
rect 71116 3296 71156 4936
rect 71212 4927 71252 4936
rect 71404 4976 71444 4985
rect 71307 4724 71349 4733
rect 71307 4684 71308 4724
rect 71348 4684 71349 4724
rect 71307 4675 71349 4684
rect 71308 4590 71348 4675
rect 71404 4397 71444 4936
rect 71499 4976 71541 4985
rect 71596 4976 71636 4985
rect 71499 4936 71500 4976
rect 71540 4936 71596 4976
rect 71499 4927 71541 4936
rect 71596 4927 71636 4936
rect 71788 4976 71828 4987
rect 71788 4901 71828 4936
rect 71883 4976 71925 4985
rect 71883 4936 71884 4976
rect 71924 4936 71925 4976
rect 71883 4927 71925 4936
rect 71787 4892 71829 4901
rect 71787 4852 71788 4892
rect 71828 4852 71829 4892
rect 71787 4843 71829 4852
rect 71884 4842 71924 4927
rect 71596 4724 71636 4733
rect 71636 4684 71924 4724
rect 71596 4675 71636 4684
rect 71403 4388 71445 4397
rect 71403 4348 71404 4388
rect 71444 4348 71445 4388
rect 71403 4339 71445 4348
rect 71307 4304 71349 4313
rect 71307 4264 71308 4304
rect 71348 4264 71349 4304
rect 71307 4255 71349 4264
rect 71116 3247 71156 3256
rect 70924 3212 70964 3221
rect 70924 2900 70964 3172
rect 70924 2860 71156 2900
rect 70924 2792 70964 2801
rect 70924 1961 70964 2752
rect 71019 2708 71061 2717
rect 71019 2668 71020 2708
rect 71060 2668 71061 2708
rect 71019 2659 71061 2668
rect 71020 2381 71060 2659
rect 71116 2624 71156 2860
rect 71211 2876 71253 2885
rect 71211 2836 71212 2876
rect 71252 2836 71253 2876
rect 71211 2827 71253 2836
rect 71116 2575 71156 2584
rect 71212 2624 71252 2827
rect 71308 2717 71348 4255
rect 71884 4136 71924 4684
rect 71884 4087 71924 4096
rect 71404 3968 71444 3977
rect 71404 3557 71444 3928
rect 71787 3716 71829 3725
rect 71787 3676 71788 3716
rect 71828 3676 71829 3716
rect 71787 3667 71829 3676
rect 71403 3548 71445 3557
rect 71595 3548 71637 3557
rect 71403 3508 71404 3548
rect 71444 3508 71445 3548
rect 71403 3499 71445 3508
rect 71500 3508 71596 3548
rect 71636 3508 71637 3548
rect 71404 3414 71444 3499
rect 71500 3464 71540 3508
rect 71595 3499 71637 3508
rect 71500 3415 71540 3424
rect 71788 3464 71828 3667
rect 71788 3415 71828 3424
rect 71691 3296 71733 3305
rect 71691 3256 71692 3296
rect 71732 3256 71733 3296
rect 71691 3247 71733 3256
rect 71692 3137 71732 3247
rect 71691 3128 71733 3137
rect 71691 3088 71692 3128
rect 71732 3088 71733 3128
rect 71691 3079 71733 3088
rect 71307 2708 71349 2717
rect 71692 2708 71732 3079
rect 71883 2792 71925 2801
rect 71883 2752 71884 2792
rect 71924 2752 71925 2792
rect 71788 2717 71828 2745
rect 71883 2743 71925 2752
rect 71787 2708 71829 2717
rect 71307 2668 71308 2708
rect 71348 2668 71349 2708
rect 71307 2659 71349 2668
rect 71691 2661 71732 2708
rect 71212 2575 71252 2584
rect 71404 2624 71444 2633
rect 71596 2624 71636 2633
rect 71444 2584 71596 2624
rect 71691 2621 71692 2661
rect 71780 2668 71788 2708
rect 71828 2668 71829 2708
rect 71780 2666 71829 2668
rect 71780 2626 71788 2666
rect 71828 2659 71829 2666
rect 71692 2612 71732 2621
rect 71788 2617 71828 2626
rect 71884 2624 71924 2743
rect 71404 2575 71444 2584
rect 71596 2575 71636 2584
rect 71884 2575 71924 2584
rect 71308 2456 71348 2465
rect 71019 2372 71061 2381
rect 71019 2332 71020 2372
rect 71060 2332 71061 2372
rect 71019 2323 71061 2332
rect 71211 2372 71253 2381
rect 71211 2332 71212 2372
rect 71252 2332 71253 2372
rect 71211 2323 71253 2332
rect 71212 2120 71252 2323
rect 71212 2071 71252 2080
rect 71308 2036 71348 2416
rect 71404 2036 71444 2045
rect 71308 1996 71404 2036
rect 71404 1987 71444 1996
rect 70923 1952 70965 1961
rect 70923 1912 70924 1952
rect 70964 1912 70965 1952
rect 70923 1903 70965 1912
rect 71787 1952 71829 1961
rect 71787 1912 71788 1952
rect 71828 1912 71829 1952
rect 71787 1903 71829 1912
rect 70827 1868 70869 1877
rect 70827 1828 70828 1868
rect 70868 1828 70869 1868
rect 70827 1819 70869 1828
rect 71788 1818 71828 1903
rect 70156 1364 70196 1373
rect 70060 1324 70156 1364
rect 70156 1315 70196 1324
rect 71884 1364 71924 1373
rect 71980 1364 72020 5608
rect 72076 4313 72116 7624
rect 72460 7328 72500 7337
rect 72364 7288 72460 7328
rect 72364 6488 72404 7288
rect 72460 7279 72500 7288
rect 72364 6439 72404 6448
rect 72171 5732 72213 5741
rect 72171 5692 72172 5732
rect 72212 5692 72213 5732
rect 72171 5683 72213 5692
rect 72172 5648 72212 5683
rect 72172 5597 72212 5608
rect 72364 5648 72404 5657
rect 72556 5648 72596 9379
rect 72940 8672 72980 10135
rect 72651 7160 72693 7169
rect 72651 7120 72652 7160
rect 72692 7120 72693 7160
rect 72651 7111 72693 7120
rect 72652 5900 72692 7111
rect 72940 6497 72980 8632
rect 72939 6488 72981 6497
rect 72939 6448 72940 6488
rect 72980 6448 72981 6488
rect 72939 6439 72981 6448
rect 72652 5851 72692 5860
rect 72404 5608 72500 5648
rect 72364 5599 72404 5608
rect 72267 5564 72309 5573
rect 72267 5524 72268 5564
rect 72308 5524 72309 5564
rect 72267 5515 72309 5524
rect 72268 5430 72308 5515
rect 72171 4976 72213 4985
rect 72171 4936 72172 4976
rect 72212 4936 72213 4976
rect 72171 4927 72213 4936
rect 72075 4304 72117 4313
rect 72075 4264 72076 4304
rect 72116 4264 72117 4304
rect 72075 4255 72117 4264
rect 72075 3632 72117 3641
rect 72075 3592 72076 3632
rect 72116 3592 72117 3632
rect 72075 3583 72117 3592
rect 72076 3464 72116 3583
rect 72172 3548 72212 4927
rect 72364 4808 72404 4817
rect 72268 4136 72308 4145
rect 72364 4136 72404 4768
rect 72460 4397 72500 5608
rect 72556 5599 72596 5608
rect 72747 5648 72789 5657
rect 72747 5608 72748 5648
rect 72788 5608 72789 5648
rect 72747 5599 72789 5608
rect 72748 5514 72788 5599
rect 73036 5396 73076 12907
rect 73324 12713 73364 16192
rect 73516 16192 73708 16232
rect 73748 16192 73940 16232
rect 73996 17032 74095 17072
rect 74188 17116 74385 17156
rect 73420 14037 73460 14046
rect 73420 13219 73460 13997
rect 73420 12965 73460 13179
rect 73419 12956 73461 12965
rect 73419 12916 73420 12956
rect 73460 12916 73461 12956
rect 73419 12907 73461 12916
rect 73323 12704 73365 12713
rect 73323 12664 73324 12704
rect 73364 12664 73365 12704
rect 73323 12655 73365 12664
rect 73516 10445 73556 16192
rect 73708 16183 73748 16192
rect 73804 16064 73844 16073
rect 73996 16064 74036 17032
rect 74188 16232 74228 17116
rect 74455 17072 74495 17472
rect 74745 17072 74785 17472
rect 74284 17032 74495 17072
rect 74572 17032 74785 17072
rect 74855 17072 74895 17472
rect 75145 17156 75185 17472
rect 74956 17116 75185 17156
rect 74855 17032 74900 17072
rect 74284 16484 74324 17032
rect 74284 16435 74324 16444
rect 74572 16232 74612 17032
rect 74668 16484 74708 16493
rect 74860 16484 74900 17032
rect 74708 16444 74900 16484
rect 74668 16435 74708 16444
rect 74228 16192 74516 16232
rect 74188 16183 74228 16192
rect 73844 16024 74036 16064
rect 73804 16015 73844 16024
rect 74283 15476 74325 15485
rect 74283 15436 74284 15476
rect 74324 15436 74325 15476
rect 74283 15427 74325 15436
rect 73803 15308 73845 15317
rect 73803 15268 73804 15308
rect 73844 15268 73845 15308
rect 73803 15259 73845 15268
rect 73611 14888 73653 14897
rect 73611 14848 73612 14888
rect 73652 14848 73653 14888
rect 73611 14839 73653 14848
rect 73612 14720 73652 14839
rect 73612 14671 73652 14680
rect 73804 14720 73844 15259
rect 74091 14888 74133 14897
rect 74091 14848 74092 14888
rect 74132 14848 74133 14888
rect 74091 14839 74133 14848
rect 73804 14671 73844 14680
rect 73900 14720 73940 14729
rect 73707 14552 73749 14561
rect 73707 14512 73708 14552
rect 73748 14512 73749 14552
rect 73707 14503 73749 14512
rect 73611 14468 73653 14477
rect 73611 14428 73612 14468
rect 73652 14428 73653 14468
rect 73611 14419 73653 14428
rect 73515 10436 73557 10445
rect 73515 10396 73516 10436
rect 73556 10396 73557 10436
rect 73515 10387 73557 10396
rect 73419 10100 73461 10109
rect 73419 10060 73420 10100
rect 73460 10060 73461 10100
rect 73419 10051 73461 10060
rect 73420 9966 73460 10051
rect 73515 8000 73557 8009
rect 73515 7960 73516 8000
rect 73556 7960 73557 8000
rect 73515 7951 73557 7960
rect 73516 7866 73556 7951
rect 73612 6656 73652 14419
rect 73708 14418 73748 14503
rect 73900 13721 73940 14680
rect 74092 14720 74132 14839
rect 74092 14671 74132 14680
rect 74188 14720 74228 14729
rect 74188 14393 74228 14680
rect 74284 14720 74324 15427
rect 74284 14671 74324 14680
rect 74380 14720 74420 14729
rect 74380 14645 74420 14680
rect 74379 14636 74421 14645
rect 74379 14596 74380 14636
rect 74420 14596 74421 14636
rect 74379 14587 74421 14596
rect 74380 14393 74420 14587
rect 74187 14384 74229 14393
rect 74187 14344 74188 14384
rect 74228 14344 74229 14384
rect 74187 14335 74229 14344
rect 74379 14384 74421 14393
rect 74379 14344 74380 14384
rect 74420 14344 74421 14384
rect 74379 14335 74421 14344
rect 74476 14132 74516 16192
rect 74092 14092 74516 14132
rect 73899 13712 73941 13721
rect 73899 13672 73900 13712
rect 73940 13672 73941 13712
rect 73899 13663 73941 13672
rect 73707 12956 73749 12965
rect 73707 12916 73708 12956
rect 73748 12916 73749 12956
rect 73707 12907 73749 12916
rect 73708 11696 73748 12907
rect 73995 12620 74037 12629
rect 73995 12580 73996 12620
rect 74036 12580 74037 12620
rect 73995 12571 74037 12580
rect 73996 11789 74036 12571
rect 73995 11780 74037 11789
rect 73995 11740 73996 11780
rect 74036 11740 74037 11780
rect 73995 11731 74037 11740
rect 73708 11647 73748 11656
rect 73804 10184 73844 10193
rect 73844 10144 73940 10184
rect 73804 10135 73844 10144
rect 73900 9344 73940 10144
rect 74092 9521 74132 14092
rect 74572 13964 74612 16192
rect 74859 16232 74901 16241
rect 74859 16192 74860 16232
rect 74900 16192 74901 16232
rect 74859 16183 74901 16192
rect 74956 16232 74996 17116
rect 75255 17072 75295 17472
rect 75545 17156 75585 17472
rect 75052 17032 75295 17072
rect 75340 17116 75585 17156
rect 75052 16484 75092 17032
rect 75052 16435 75092 16444
rect 75340 16241 75380 17116
rect 75655 17072 75695 17472
rect 75945 17249 75985 17472
rect 75944 17240 75986 17249
rect 75944 17200 75945 17240
rect 75985 17200 75986 17240
rect 75944 17191 75986 17200
rect 76055 17072 76095 17472
rect 75436 17032 75695 17072
rect 75820 17032 76095 17072
rect 75436 16484 75476 17032
rect 75436 16435 75476 16444
rect 75820 16484 75860 17032
rect 76345 16988 76385 17472
rect 76455 17072 76495 17472
rect 76455 17032 76532 17072
rect 76345 16948 76436 16988
rect 75820 16435 75860 16444
rect 74667 15392 74709 15401
rect 74667 15352 74668 15392
rect 74708 15352 74709 15392
rect 74667 15343 74709 15352
rect 74668 14720 74708 15343
rect 74763 14804 74805 14813
rect 74763 14764 74764 14804
rect 74804 14764 74805 14804
rect 74763 14755 74805 14764
rect 74668 14671 74708 14680
rect 74667 14048 74709 14057
rect 74667 14008 74668 14048
rect 74708 14008 74709 14048
rect 74667 13999 74709 14008
rect 74764 14048 74804 14755
rect 74860 14477 74900 16183
rect 74956 16157 74996 16192
rect 75339 16232 75381 16241
rect 75339 16192 75340 16232
rect 75380 16192 75381 16232
rect 75339 16183 75381 16192
rect 75723 16232 75765 16241
rect 75723 16192 75724 16232
rect 75764 16192 75765 16232
rect 76396 16232 76436 16948
rect 76492 16484 76532 17032
rect 76745 16988 76785 17472
rect 76855 17072 76895 17472
rect 77145 17072 77185 17472
rect 77255 17072 77295 17472
rect 77545 17156 77585 17472
rect 77452 17116 77585 17156
rect 76855 17032 76916 17072
rect 77145 17032 77204 17072
rect 77255 17032 77300 17072
rect 76745 16948 76820 16988
rect 76492 16435 76532 16444
rect 76588 16232 76628 16241
rect 76396 16192 76588 16232
rect 76780 16232 76820 16948
rect 76876 16484 76916 17032
rect 76876 16435 76916 16444
rect 77164 16241 77204 17032
rect 77260 16484 77300 17032
rect 77260 16435 77300 16444
rect 76972 16232 77012 16241
rect 76780 16192 76972 16232
rect 75723 16183 75765 16192
rect 74955 16148 74997 16157
rect 74955 16108 74956 16148
rect 74996 16108 74997 16148
rect 74955 16099 74997 16108
rect 74956 16068 74996 16099
rect 75340 16098 75380 16183
rect 75724 16098 75764 16183
rect 76588 16073 76628 16192
rect 76587 16064 76629 16073
rect 76587 16024 76588 16064
rect 76628 16024 76629 16064
rect 76587 16015 76629 16024
rect 76972 15821 77012 16192
rect 77163 16232 77205 16241
rect 77452 16232 77492 17116
rect 77655 17072 77695 17472
rect 77945 17156 77985 17472
rect 77548 17032 77695 17072
rect 77836 17116 77985 17156
rect 77548 16484 77588 17032
rect 77548 16435 77588 16444
rect 77163 16192 77164 16232
rect 77204 16192 77205 16232
rect 77163 16183 77205 16192
rect 77356 16192 77452 16232
rect 77164 16098 77204 16183
rect 76971 15812 77013 15821
rect 76971 15772 76972 15812
rect 77012 15772 77013 15812
rect 76971 15763 77013 15772
rect 75147 15560 75189 15569
rect 75147 15520 75148 15560
rect 75188 15520 75189 15560
rect 75147 15511 75189 15520
rect 75340 15560 75380 15569
rect 75380 15520 75572 15560
rect 75340 15511 75380 15520
rect 75148 15426 75188 15511
rect 75244 15317 75284 15402
rect 75243 15308 75285 15317
rect 75243 15268 75244 15308
rect 75284 15268 75285 15308
rect 75243 15259 75285 15268
rect 75112 15140 75480 15149
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75112 15091 75480 15100
rect 75340 14972 75380 14981
rect 75532 14972 75572 15520
rect 76684 15392 76724 15401
rect 75627 15308 75669 15317
rect 75627 15268 75628 15308
rect 75668 15268 75669 15308
rect 75627 15259 75669 15268
rect 75380 14932 75572 14972
rect 75340 14923 75380 14932
rect 75628 14897 75668 15259
rect 75627 14888 75669 14897
rect 75627 14848 75628 14888
rect 75668 14848 75669 14888
rect 75627 14839 75669 14848
rect 75724 14848 76244 14888
rect 74956 14720 74996 14729
rect 74956 14561 74996 14680
rect 75627 14720 75669 14729
rect 75627 14680 75628 14720
rect 75668 14680 75669 14720
rect 75627 14671 75669 14680
rect 75051 14636 75093 14645
rect 75051 14596 75052 14636
rect 75092 14596 75093 14636
rect 75051 14587 75093 14596
rect 74955 14552 74997 14561
rect 74955 14512 74956 14552
rect 74996 14512 74997 14552
rect 74955 14503 74997 14512
rect 75052 14502 75092 14587
rect 75628 14586 75668 14671
rect 75724 14636 75764 14848
rect 75819 14720 75861 14729
rect 75819 14680 75820 14720
rect 75860 14680 75861 14720
rect 75819 14671 75861 14680
rect 75916 14720 75956 14729
rect 75724 14587 75764 14596
rect 75820 14586 75860 14671
rect 74859 14468 74901 14477
rect 74859 14428 74860 14468
rect 74900 14428 74901 14468
rect 74859 14419 74901 14428
rect 75916 14132 75956 14680
rect 76204 14720 76244 14848
rect 76204 14671 76244 14680
rect 76588 14720 76628 14729
rect 76684 14720 76724 15352
rect 76628 14680 76724 14720
rect 76588 14671 76628 14680
rect 76011 14552 76053 14561
rect 76011 14512 76012 14552
rect 76052 14512 76053 14552
rect 77356 14552 77396 16192
rect 77452 16183 77492 16192
rect 77836 16232 77876 17116
rect 78055 17072 78095 17472
rect 78345 17156 78385 17472
rect 77932 17032 78095 17072
rect 78220 17116 78385 17156
rect 77932 16484 77972 17032
rect 77932 16435 77972 16444
rect 78220 16232 78260 17116
rect 78455 17072 78495 17472
rect 78745 17156 78785 17472
rect 78316 17032 78495 17072
rect 78604 17116 78785 17156
rect 78316 16484 78356 17032
rect 78316 16435 78356 16444
rect 78604 16232 78644 17116
rect 78855 17072 78895 17472
rect 78987 17156 79029 17165
rect 78987 17116 78988 17156
rect 79028 17116 79029 17156
rect 78987 17107 79029 17116
rect 78700 17032 78895 17072
rect 78700 16484 78740 17032
rect 78700 16435 78740 16444
rect 78988 16484 79028 17107
rect 79145 17072 79185 17472
rect 79255 17156 79295 17472
rect 79371 17156 79413 17165
rect 79255 17116 79316 17156
rect 79145 17032 79220 17072
rect 78988 16435 79028 16444
rect 78891 16232 78933 16241
rect 77876 16192 77972 16232
rect 77836 16183 77876 16192
rect 77452 14720 77492 14729
rect 77492 14680 77684 14720
rect 77452 14671 77492 14680
rect 77356 14512 77588 14552
rect 76011 14503 76053 14512
rect 75916 14083 75956 14092
rect 74764 13999 74804 14008
rect 74956 14048 74996 14059
rect 74188 13924 74612 13964
rect 74091 9512 74133 9521
rect 74091 9472 74092 9512
rect 74132 9472 74133 9512
rect 74091 9463 74133 9472
rect 73900 9295 73940 9304
rect 74092 8924 74132 9463
rect 74188 9008 74228 13924
rect 74572 13796 74612 13805
rect 74668 13796 74708 13999
rect 74956 13973 74996 14008
rect 75052 14048 75092 14057
rect 74955 13964 74997 13973
rect 74955 13924 74956 13964
rect 74996 13924 74997 13964
rect 74955 13915 74997 13924
rect 74859 13880 74901 13889
rect 74859 13840 74860 13880
rect 74900 13840 74901 13880
rect 74859 13831 74901 13840
rect 74612 13756 74708 13796
rect 74764 13796 74804 13807
rect 74572 13747 74612 13756
rect 74764 13721 74804 13756
rect 74763 13712 74805 13721
rect 74763 13672 74764 13712
rect 74804 13672 74805 13712
rect 74763 13663 74805 13672
rect 74860 13553 74900 13831
rect 75052 13796 75092 14008
rect 75820 14048 75860 14057
rect 75820 13805 75860 14008
rect 76012 14048 76052 14503
rect 76352 14384 76720 14393
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76352 14335 76720 14344
rect 77163 14216 77205 14225
rect 77163 14176 77164 14216
rect 77204 14176 77205 14216
rect 77163 14167 77205 14176
rect 76972 14048 77012 14057
rect 76012 13999 76052 14008
rect 76492 14008 76972 14048
rect 74956 13756 75092 13796
rect 75819 13796 75861 13805
rect 75819 13756 75820 13796
rect 75860 13756 75861 13796
rect 74859 13544 74901 13553
rect 74859 13504 74860 13544
rect 74900 13504 74901 13544
rect 74859 13495 74901 13504
rect 74572 13385 74612 13470
rect 74956 13385 74996 13756
rect 75819 13747 75861 13756
rect 75112 13628 75480 13637
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75112 13579 75480 13588
rect 75147 13460 75189 13469
rect 75147 13420 75148 13460
rect 75188 13420 75189 13460
rect 75147 13411 75189 13420
rect 76492 13460 76532 14008
rect 76972 13999 77012 14008
rect 76492 13411 76532 13420
rect 74379 13376 74421 13385
rect 74379 13336 74380 13376
rect 74420 13336 74421 13376
rect 74379 13327 74421 13336
rect 74571 13376 74613 13385
rect 74571 13336 74572 13376
rect 74612 13336 74613 13376
rect 74571 13327 74613 13336
rect 74955 13376 74997 13385
rect 74955 13336 74956 13376
rect 74996 13336 74997 13376
rect 74955 13327 74997 13336
rect 74283 13208 74325 13217
rect 74283 13168 74284 13208
rect 74324 13168 74325 13208
rect 74283 13159 74325 13168
rect 74284 12536 74324 13159
rect 74380 12704 74420 13327
rect 74763 13208 74805 13217
rect 74763 13168 74764 13208
rect 74804 13168 74805 13208
rect 74763 13159 74805 13168
rect 74860 13208 74900 13217
rect 74764 13074 74804 13159
rect 74860 12980 74900 13168
rect 74956 13208 74996 13219
rect 74956 13133 74996 13168
rect 75051 13208 75093 13217
rect 75051 13168 75052 13208
rect 75092 13168 75093 13208
rect 75051 13159 75093 13168
rect 74955 13124 74997 13133
rect 74955 13084 74956 13124
rect 74996 13084 74997 13124
rect 74955 13075 74997 13084
rect 75052 13074 75092 13159
rect 75148 13133 75188 13411
rect 76108 13376 76148 13385
rect 77068 13376 77108 13385
rect 75723 13292 75765 13301
rect 75723 13252 75724 13292
rect 75764 13252 75765 13292
rect 75723 13243 75765 13252
rect 75436 13208 75476 13217
rect 75147 13124 75189 13133
rect 75147 13084 75148 13124
rect 75188 13084 75189 13124
rect 75147 13075 75189 13084
rect 75148 12980 75188 13075
rect 75436 13040 75476 13168
rect 75724 13208 75764 13243
rect 75724 13157 75764 13168
rect 75819 13208 75861 13217
rect 75819 13168 75820 13208
rect 75860 13168 75861 13208
rect 75819 13159 75861 13168
rect 75820 13074 75860 13159
rect 75531 13040 75573 13049
rect 75436 13000 75532 13040
rect 75572 13000 75573 13040
rect 75531 12991 75573 13000
rect 74668 12940 74900 12980
rect 74956 12940 75188 12980
rect 74380 12655 74420 12664
rect 74475 12704 74517 12713
rect 74475 12664 74476 12704
rect 74516 12664 74517 12704
rect 74475 12655 74517 12664
rect 74284 12487 74324 12496
rect 74476 12536 74516 12655
rect 74476 12487 74516 12496
rect 74572 12536 74612 12545
rect 74572 12377 74612 12496
rect 74571 12368 74613 12377
rect 74571 12328 74572 12368
rect 74612 12328 74613 12368
rect 74571 12319 74613 12328
rect 74668 12200 74708 12940
rect 74764 12629 74804 12673
rect 74763 12620 74805 12629
rect 74763 12580 74764 12620
rect 74804 12580 74805 12620
rect 74763 12578 74805 12580
rect 74763 12571 74764 12578
rect 74804 12571 74805 12578
rect 74764 12529 74804 12538
rect 74956 12536 74996 12940
rect 74956 12487 74996 12496
rect 75052 12536 75092 12545
rect 74764 12377 74804 12462
rect 74763 12368 74805 12377
rect 74763 12328 74764 12368
rect 74804 12328 74805 12368
rect 74763 12319 74805 12328
rect 75052 12284 75092 12496
rect 74956 12244 75092 12284
rect 74668 12160 74804 12200
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 74764 11024 74804 12160
rect 74956 11957 74996 12244
rect 75112 12116 75480 12125
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75112 12067 75480 12076
rect 74860 11948 74900 11957
rect 74955 11948 74997 11957
rect 74900 11908 74956 11948
rect 74996 11908 74997 11948
rect 74860 11899 74900 11908
rect 74955 11899 74997 11908
rect 74859 11360 74901 11369
rect 74859 11320 74860 11360
rect 74900 11320 74901 11360
rect 74859 11311 74901 11320
rect 74668 10890 74708 10975
rect 74764 10352 74804 10984
rect 74572 10312 74804 10352
rect 74860 11024 74900 11311
rect 74572 9605 74612 10312
rect 74667 10184 74709 10193
rect 74667 10144 74668 10184
rect 74708 10144 74804 10184
rect 74667 10135 74709 10144
rect 74668 10050 74708 10135
rect 74571 9596 74613 9605
rect 74571 9556 74572 9596
rect 74612 9556 74613 9596
rect 74571 9547 74613 9556
rect 74188 8968 74420 9008
rect 74092 8875 74132 8884
rect 74284 8840 74324 8849
rect 73900 8000 73940 8009
rect 74284 8000 74324 8800
rect 73940 7960 74324 8000
rect 73900 7951 73940 7960
rect 74380 6656 74420 8968
rect 74764 8000 74804 10144
rect 74860 9689 74900 10984
rect 74956 11024 74996 11899
rect 75340 11696 75380 11705
rect 75340 11528 75380 11656
rect 75435 11528 75477 11537
rect 75532 11528 75572 12991
rect 76108 12980 76148 13336
rect 76780 13336 77068 13376
rect 76491 13208 76533 13217
rect 76491 13168 76492 13208
rect 76532 13168 76533 13208
rect 76491 13159 76533 13168
rect 76684 13208 76724 13217
rect 76492 13074 76532 13159
rect 76684 12980 76724 13168
rect 76780 13208 76820 13336
rect 77068 13327 77108 13336
rect 77164 13301 77204 14167
rect 77356 14048 77396 14057
rect 77356 13376 77396 14008
rect 77452 13376 77492 13385
rect 77356 13336 77452 13376
rect 77452 13327 77492 13336
rect 77163 13292 77205 13301
rect 77163 13252 77164 13292
rect 77204 13252 77205 13292
rect 77163 13243 77205 13252
rect 76780 13159 76820 13168
rect 76972 13208 77012 13219
rect 76972 13133 77012 13168
rect 77164 13208 77204 13243
rect 77164 13158 77204 13168
rect 76971 13124 77013 13133
rect 76971 13084 76972 13124
rect 77012 13084 77013 13124
rect 76971 13075 77013 13084
rect 76108 12940 76244 12980
rect 76684 12940 76820 12980
rect 76107 12704 76149 12713
rect 76107 12664 76108 12704
rect 76148 12664 76149 12704
rect 76107 12655 76149 12664
rect 75819 12620 75861 12629
rect 75819 12580 75820 12620
rect 75860 12580 75861 12620
rect 75819 12571 75861 12580
rect 76108 12620 76148 12655
rect 75723 11948 75765 11957
rect 75723 11908 75724 11948
rect 75764 11908 75765 11948
rect 75723 11899 75765 11908
rect 75628 11705 75668 11790
rect 75627 11696 75669 11705
rect 75627 11656 75628 11696
rect 75668 11656 75669 11696
rect 75627 11647 75669 11656
rect 75724 11696 75764 11899
rect 75724 11647 75764 11656
rect 75820 11528 75860 12571
rect 76108 12569 76148 12580
rect 76012 12536 76052 12545
rect 76012 12032 76052 12496
rect 76204 12536 76244 12940
rect 76352 12872 76720 12881
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76352 12823 76720 12832
rect 76780 12713 76820 12940
rect 76779 12704 76821 12713
rect 76779 12664 76780 12704
rect 76820 12664 76821 12704
rect 76779 12655 76821 12664
rect 76876 12545 76916 12630
rect 76204 12487 76244 12496
rect 76395 12536 76437 12545
rect 76395 12496 76396 12536
rect 76436 12496 76437 12536
rect 76395 12487 76437 12496
rect 76875 12536 76917 12545
rect 76875 12496 76876 12536
rect 76916 12496 76917 12536
rect 76875 12487 76917 12496
rect 76012 11992 76340 12032
rect 76012 11864 76052 11873
rect 76052 11824 76148 11864
rect 76012 11815 76052 11824
rect 75340 11488 75436 11528
rect 75476 11488 75572 11528
rect 75724 11488 75860 11528
rect 76011 11528 76053 11537
rect 76011 11488 76012 11528
rect 76052 11488 76053 11528
rect 75435 11479 75477 11488
rect 75339 11360 75381 11369
rect 75339 11320 75340 11360
rect 75380 11320 75381 11360
rect 75339 11311 75381 11320
rect 75243 11192 75285 11201
rect 75243 11152 75244 11192
rect 75284 11152 75285 11192
rect 75243 11143 75285 11152
rect 75244 11058 75284 11143
rect 74956 10975 74996 10984
rect 75147 11024 75189 11033
rect 75147 10984 75148 11024
rect 75188 10984 75189 11024
rect 75147 10975 75189 10984
rect 75340 11024 75380 11311
rect 75340 10975 75380 10984
rect 75436 11024 75476 11033
rect 75148 10890 75188 10975
rect 75436 10856 75476 10984
rect 75628 11024 75668 11033
rect 75724 11024 75764 11488
rect 76011 11479 76053 11488
rect 75668 10984 75764 11024
rect 75628 10975 75668 10984
rect 75628 10856 75668 10865
rect 75436 10816 75628 10856
rect 75628 10807 75668 10816
rect 75112 10604 75480 10613
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75112 10555 75480 10564
rect 75724 10268 75764 10984
rect 75819 11024 75861 11033
rect 75819 10984 75820 11024
rect 75860 10984 75861 11024
rect 75819 10975 75861 10984
rect 75916 11024 75956 11033
rect 75820 10890 75860 10975
rect 75916 10445 75956 10984
rect 75820 10436 75860 10445
rect 75915 10436 75957 10445
rect 75860 10396 75916 10436
rect 75956 10396 75957 10436
rect 75820 10387 75860 10396
rect 75915 10387 75957 10396
rect 75916 10302 75956 10387
rect 75436 10228 75764 10268
rect 74859 9680 74901 9689
rect 74859 9640 74860 9680
rect 74900 9640 74901 9680
rect 74859 9631 74901 9640
rect 74860 8093 74900 9631
rect 75436 9512 75476 10228
rect 76012 10184 76052 11479
rect 76108 11024 76148 11824
rect 76203 11696 76245 11705
rect 76203 11656 76204 11696
rect 76244 11656 76245 11696
rect 76203 11647 76245 11656
rect 76204 11108 76244 11647
rect 76300 11537 76340 11992
rect 76396 11948 76436 12487
rect 76972 12368 77012 13075
rect 77548 12980 77588 14512
rect 77644 14057 77684 14680
rect 77643 14048 77685 14057
rect 77643 14008 77644 14048
rect 77684 14008 77685 14048
rect 77643 13999 77685 14008
rect 77452 12940 77588 12980
rect 77644 12965 77684 13999
rect 77932 12980 77972 16192
rect 78260 16192 78356 16232
rect 78220 16183 78260 16192
rect 78219 14048 78261 14057
rect 78219 14008 78220 14048
rect 78260 14008 78261 14048
rect 78219 13999 78261 14008
rect 78220 13914 78260 13999
rect 77643 12956 77685 12965
rect 76396 11899 76436 11908
rect 76876 12328 77012 12368
rect 77260 12536 77300 12545
rect 76396 11696 76436 11707
rect 76396 11621 76436 11656
rect 76587 11696 76629 11705
rect 76587 11656 76588 11696
rect 76628 11656 76629 11696
rect 76587 11647 76629 11656
rect 76684 11696 76724 11705
rect 76876 11696 76916 12328
rect 77260 11864 77300 12496
rect 77356 11864 77396 11873
rect 77260 11824 77356 11864
rect 77356 11815 77396 11824
rect 77067 11780 77109 11789
rect 77067 11740 77068 11780
rect 77108 11740 77109 11780
rect 77067 11731 77109 11740
rect 76724 11656 76820 11696
rect 76684 11647 76724 11656
rect 76395 11612 76437 11621
rect 76395 11572 76396 11612
rect 76436 11572 76437 11612
rect 76395 11563 76437 11572
rect 76588 11562 76628 11647
rect 76299 11528 76341 11537
rect 76299 11488 76300 11528
rect 76340 11488 76341 11528
rect 76780 11528 76820 11656
rect 76876 11647 76916 11656
rect 77068 11696 77108 11731
rect 77068 11645 77108 11656
rect 76972 11612 77012 11621
rect 76972 11528 77012 11572
rect 77163 11612 77205 11621
rect 77163 11572 77164 11612
rect 77204 11572 77205 11612
rect 77163 11563 77205 11572
rect 76780 11488 77012 11528
rect 76299 11479 76341 11488
rect 76352 11360 76720 11369
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76352 11311 76720 11320
rect 76299 11192 76341 11201
rect 76299 11152 76300 11192
rect 76340 11152 76341 11192
rect 76299 11143 76341 11152
rect 76204 11059 76244 11068
rect 76108 10975 76148 10984
rect 76300 11024 76340 11143
rect 77059 11037 77099 11046
rect 76204 10184 76244 10193
rect 76012 10144 76204 10184
rect 75915 10100 75957 10109
rect 75915 10060 75916 10100
rect 75956 10060 75957 10100
rect 75915 10051 75957 10060
rect 75820 10016 75860 10025
rect 75531 9848 75573 9857
rect 75531 9808 75532 9848
rect 75572 9808 75573 9848
rect 75531 9799 75573 9808
rect 75532 9680 75572 9799
rect 75532 9631 75572 9640
rect 75723 9680 75765 9689
rect 75723 9640 75724 9680
rect 75764 9640 75765 9680
rect 75723 9631 75765 9640
rect 75627 9596 75669 9605
rect 75627 9556 75628 9596
rect 75668 9556 75669 9596
rect 75627 9547 75669 9556
rect 75628 9512 75668 9547
rect 75436 9472 75572 9512
rect 75112 9092 75480 9101
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75112 9043 75480 9052
rect 75532 8672 75572 9472
rect 75724 9533 75764 9631
rect 75724 9484 75764 9493
rect 75820 9533 75860 9976
rect 75820 9484 75860 9493
rect 75628 9461 75668 9472
rect 75916 9344 75956 10051
rect 76011 9848 76053 9857
rect 76011 9808 76012 9848
rect 76052 9808 76053 9848
rect 76011 9799 76053 9808
rect 76012 9512 76052 9799
rect 76108 9596 76148 10144
rect 76204 10135 76244 10144
rect 76300 10109 76340 10984
rect 76683 11024 76725 11033
rect 76683 10984 76684 11024
rect 76724 10984 76725 11024
rect 76683 10975 76725 10984
rect 76972 10997 77059 11024
rect 76972 10984 77099 10997
rect 76492 10940 76532 10949
rect 76396 10900 76492 10940
rect 76299 10100 76341 10109
rect 76299 10060 76300 10100
rect 76340 10060 76341 10100
rect 76299 10051 76341 10060
rect 76396 10025 76436 10900
rect 76492 10891 76532 10900
rect 76684 10772 76724 10975
rect 76724 10732 76820 10772
rect 76684 10723 76724 10732
rect 76587 10436 76629 10445
rect 76587 10396 76588 10436
rect 76628 10396 76629 10436
rect 76587 10387 76629 10396
rect 76491 10268 76533 10277
rect 76491 10228 76492 10268
rect 76532 10228 76533 10268
rect 76491 10219 76533 10228
rect 76492 10184 76532 10219
rect 76492 10133 76532 10144
rect 76588 10184 76628 10387
rect 76588 10135 76628 10144
rect 76395 10016 76437 10025
rect 76395 9976 76396 10016
rect 76436 9976 76437 10016
rect 76395 9967 76437 9976
rect 76352 9848 76720 9857
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76352 9799 76720 9808
rect 76491 9680 76533 9689
rect 76491 9640 76492 9680
rect 76532 9640 76533 9680
rect 76491 9631 76533 9640
rect 76107 9556 76148 9596
rect 76107 9512 76147 9556
rect 76204 9525 76244 9607
rect 76107 9472 76148 9512
rect 76012 9463 76052 9472
rect 76012 9344 76052 9353
rect 75916 9304 76012 9344
rect 76012 9295 76052 9304
rect 75819 9260 75861 9269
rect 75819 9220 75820 9260
rect 75860 9220 75861 9260
rect 75819 9211 75861 9220
rect 75628 8672 75668 8681
rect 75532 8632 75628 8672
rect 75628 8336 75668 8632
rect 75820 8672 75860 9211
rect 76108 9176 76148 9472
rect 76203 9472 76204 9521
rect 76244 9472 76245 9521
rect 76203 9463 76245 9472
rect 76300 9512 76340 9521
rect 76108 9136 76244 9176
rect 75723 8588 75765 8597
rect 75723 8548 75724 8588
rect 75764 8548 75765 8588
rect 75723 8539 75765 8548
rect 75724 8454 75764 8539
rect 75628 8296 75764 8336
rect 74859 8084 74901 8093
rect 74859 8044 74860 8084
rect 74900 8044 74901 8084
rect 74859 8035 74901 8044
rect 74764 7951 74804 7960
rect 73612 6616 73748 6656
rect 73227 6488 73269 6497
rect 73227 6448 73228 6488
rect 73268 6448 73269 6488
rect 73227 6439 73269 6448
rect 73611 6488 73653 6497
rect 73611 6448 73612 6488
rect 73652 6448 73653 6488
rect 73611 6439 73653 6448
rect 73228 6354 73268 6439
rect 73612 5900 73652 6439
rect 73612 5851 73652 5860
rect 72652 5356 73076 5396
rect 72459 4388 72501 4397
rect 72459 4348 72460 4388
rect 72500 4348 72501 4388
rect 72459 4339 72501 4348
rect 72308 4096 72404 4136
rect 72268 4087 72308 4096
rect 72172 3499 72212 3508
rect 72267 3548 72309 3557
rect 72267 3508 72268 3548
rect 72308 3508 72309 3548
rect 72267 3499 72309 3508
rect 72076 3415 72116 3424
rect 72268 3464 72308 3499
rect 72268 3413 72308 3424
rect 72459 3464 72501 3473
rect 72459 3424 72460 3464
rect 72500 3424 72501 3464
rect 72459 3415 72501 3424
rect 72460 3330 72500 3415
rect 72652 2876 72692 5356
rect 72843 4388 72885 4397
rect 72843 4348 72844 4388
rect 72884 4348 72885 4388
rect 72843 4339 72885 4348
rect 72747 3464 72789 3473
rect 72747 3424 72748 3464
rect 72788 3424 72789 3464
rect 72747 3415 72789 3424
rect 72844 3464 72884 4339
rect 73708 4313 73748 6616
rect 74380 6607 74420 6616
rect 74860 6581 74900 8035
rect 75531 8000 75573 8009
rect 75531 7960 75532 8000
rect 75572 7960 75573 8000
rect 75531 7951 75573 7960
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 75532 7412 75572 7951
rect 75627 7916 75669 7925
rect 75627 7876 75628 7916
rect 75668 7876 75669 7916
rect 75627 7867 75669 7876
rect 75532 7363 75572 7372
rect 75435 7244 75477 7253
rect 75435 7204 75436 7244
rect 75476 7204 75477 7244
rect 75435 7195 75477 7204
rect 75436 6992 75476 7195
rect 75532 7160 75572 7169
rect 75628 7160 75668 7867
rect 75724 7841 75764 8296
rect 75723 7832 75765 7841
rect 75723 7792 75724 7832
rect 75764 7792 75765 7832
rect 75723 7783 75765 7792
rect 75820 7337 75860 8632
rect 75916 8672 75956 8681
rect 75916 8513 75956 8632
rect 76204 8672 76244 9136
rect 76204 8588 76244 8632
rect 76300 8597 76340 9472
rect 76492 9428 76532 9631
rect 76587 9596 76629 9605
rect 76587 9556 76588 9596
rect 76628 9556 76629 9596
rect 76587 9547 76629 9556
rect 76492 9379 76532 9388
rect 76588 9260 76628 9547
rect 76780 9437 76820 10732
rect 76876 10436 76916 10445
rect 76972 10436 77012 10984
rect 77164 10940 77204 11563
rect 77259 11192 77301 11201
rect 77259 11152 77260 11192
rect 77300 11152 77301 11192
rect 77259 11143 77301 11152
rect 77260 11024 77300 11143
rect 77260 10975 77300 10984
rect 76916 10396 77012 10436
rect 77068 10900 77204 10940
rect 76876 10387 76916 10396
rect 77068 10352 77108 10900
rect 77164 10772 77204 10781
rect 77204 10732 77300 10772
rect 77164 10723 77204 10732
rect 76972 10312 77108 10352
rect 76875 10100 76917 10109
rect 76875 10060 76876 10100
rect 76916 10060 76917 10100
rect 76875 10051 76917 10060
rect 76779 9428 76821 9437
rect 76779 9388 76780 9428
rect 76820 9388 76821 9428
rect 76779 9379 76821 9388
rect 76492 9220 76628 9260
rect 76683 9260 76725 9269
rect 76683 9220 76684 9260
rect 76724 9220 76725 9260
rect 76492 8672 76532 9220
rect 76683 9211 76725 9220
rect 76684 9126 76724 9211
rect 76876 9008 76916 10051
rect 76492 8623 76532 8632
rect 76780 8968 76916 9008
rect 76972 9512 77012 10312
rect 77068 10100 77108 10109
rect 77068 9680 77108 10060
rect 77164 9680 77204 9689
rect 77068 9640 77164 9680
rect 77164 9631 77204 9640
rect 77260 9521 77300 10732
rect 77452 10352 77492 12940
rect 77643 12916 77644 12956
rect 77684 12916 77685 12956
rect 77643 12907 77685 12916
rect 77740 12940 77972 12980
rect 77644 12545 77684 12907
rect 77643 12536 77685 12545
rect 77643 12496 77644 12536
rect 77684 12496 77685 12536
rect 77643 12487 77685 12496
rect 77356 10312 77492 10352
rect 77644 10856 77684 10865
rect 77356 9689 77396 10312
rect 77452 10184 77492 10193
rect 77644 10184 77684 10816
rect 77740 10277 77780 12940
rect 78123 12536 78165 12545
rect 78123 12496 78124 12536
rect 78164 12496 78165 12536
rect 78123 12487 78165 12496
rect 78124 12402 78164 12487
rect 78316 12293 78356 16192
rect 78644 16192 78740 16232
rect 78604 16183 78644 16192
rect 78411 15812 78453 15821
rect 78411 15772 78412 15812
rect 78452 15772 78453 15812
rect 78411 15763 78453 15772
rect 78315 12284 78357 12293
rect 78315 12244 78316 12284
rect 78356 12244 78357 12284
rect 78315 12235 78357 12244
rect 78316 11789 78356 12235
rect 78315 11780 78357 11789
rect 78315 11740 78316 11780
rect 78356 11740 78357 11780
rect 78315 11731 78357 11740
rect 77739 10268 77781 10277
rect 77739 10228 77740 10268
rect 77780 10228 77781 10268
rect 77739 10219 77781 10228
rect 77492 10144 77684 10184
rect 77452 10135 77492 10144
rect 77355 9680 77397 9689
rect 77355 9640 77356 9680
rect 77396 9640 77397 9680
rect 77355 9631 77397 9640
rect 77548 9521 77588 9606
rect 77068 9512 77108 9521
rect 76972 9472 77068 9512
rect 76012 8548 76244 8588
rect 76299 8588 76341 8597
rect 76299 8548 76300 8588
rect 76340 8548 76341 8588
rect 75915 8504 75957 8513
rect 75915 8464 75916 8504
rect 75956 8464 75957 8504
rect 75915 8455 75957 8464
rect 75916 8177 75956 8455
rect 75915 8168 75957 8177
rect 75915 8128 75916 8168
rect 75956 8128 75957 8168
rect 75915 8119 75957 8128
rect 76012 8000 76052 8548
rect 76299 8539 76341 8548
rect 76587 8588 76629 8597
rect 76587 8548 76588 8588
rect 76628 8548 76629 8588
rect 76587 8539 76629 8548
rect 76588 8454 76628 8539
rect 76203 8420 76245 8429
rect 76203 8380 76204 8420
rect 76244 8380 76245 8420
rect 76203 8371 76245 8380
rect 76108 8009 76148 8094
rect 75916 7960 76052 8000
rect 76107 8000 76149 8009
rect 76107 7960 76108 8000
rect 76148 7960 76149 8000
rect 75819 7328 75861 7337
rect 75819 7288 75820 7328
rect 75860 7288 75861 7328
rect 75819 7279 75861 7288
rect 75572 7120 75668 7160
rect 75723 7160 75765 7169
rect 75723 7120 75724 7160
rect 75764 7120 75765 7160
rect 75532 7111 75572 7120
rect 75723 7111 75765 7120
rect 75820 7160 75860 7171
rect 75724 7026 75764 7111
rect 75820 7085 75860 7120
rect 75819 7076 75861 7085
rect 75819 7036 75820 7076
rect 75860 7036 75861 7076
rect 75916 7076 75956 7960
rect 76107 7951 76149 7960
rect 76204 8000 76244 8371
rect 76352 8336 76720 8345
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76352 8287 76720 8296
rect 76395 8168 76437 8177
rect 76780 8168 76820 8968
rect 76395 8128 76396 8168
rect 76436 8128 76437 8168
rect 76395 8119 76437 8128
rect 76588 8128 76820 8168
rect 76876 8840 76916 8849
rect 76299 8084 76341 8093
rect 76299 8044 76300 8084
rect 76340 8044 76341 8084
rect 76299 8035 76341 8044
rect 76011 7832 76053 7841
rect 76011 7792 76012 7832
rect 76052 7792 76053 7832
rect 76011 7783 76053 7792
rect 76012 7171 76052 7783
rect 76204 7421 76244 7960
rect 76300 8000 76340 8035
rect 76300 7949 76340 7960
rect 76396 8000 76436 8119
rect 76396 7951 76436 7960
rect 76588 8000 76628 8128
rect 76203 7412 76245 7421
rect 76203 7372 76204 7412
rect 76244 7372 76245 7412
rect 76203 7363 76245 7372
rect 76588 7253 76628 7960
rect 76780 8000 76820 8009
rect 76876 8000 76916 8800
rect 76820 7960 76916 8000
rect 76972 8000 77012 9472
rect 77068 9463 77108 9472
rect 77259 9512 77301 9521
rect 77259 9472 77260 9512
rect 77300 9472 77301 9512
rect 77259 9463 77301 9472
rect 77356 9512 77396 9521
rect 77260 9378 77300 9463
rect 77356 9344 77396 9472
rect 77547 9512 77589 9521
rect 77547 9472 77548 9512
rect 77588 9472 77589 9512
rect 77547 9463 77589 9472
rect 77740 9512 77780 10219
rect 78315 10184 78357 10193
rect 78315 10144 78316 10184
rect 78356 10144 78357 10184
rect 78315 10135 78357 10144
rect 78123 9680 78165 9689
rect 78123 9640 78124 9680
rect 78164 9640 78165 9680
rect 78123 9631 78165 9640
rect 77740 9463 77780 9472
rect 77931 9512 77973 9521
rect 77931 9472 77932 9512
rect 77972 9472 77973 9512
rect 77931 9463 77973 9472
rect 78124 9512 78164 9631
rect 78124 9463 78164 9472
rect 77932 9378 77972 9463
rect 77644 9344 77684 9353
rect 77356 9304 77644 9344
rect 77644 9295 77684 9304
rect 78028 9260 78068 9269
rect 77355 9176 77397 9185
rect 77355 9136 77356 9176
rect 77396 9136 77397 9176
rect 77355 9127 77397 9136
rect 77068 8588 77108 8597
rect 77068 8168 77108 8548
rect 77068 8119 77108 8128
rect 76780 7951 76820 7960
rect 76972 7832 77012 7960
rect 76780 7792 77012 7832
rect 77164 8000 77204 8009
rect 76684 7748 76724 7757
rect 76203 7244 76245 7253
rect 76203 7204 76204 7244
rect 76244 7204 76245 7244
rect 76203 7195 76245 7204
rect 76587 7244 76629 7253
rect 76587 7204 76588 7244
rect 76628 7204 76629 7244
rect 76587 7195 76629 7204
rect 76012 7122 76052 7131
rect 76108 7085 76148 7170
rect 76204 7160 76244 7195
rect 76684 7169 76724 7708
rect 76204 7109 76244 7120
rect 76300 7160 76340 7169
rect 76107 7076 76149 7085
rect 75916 7036 76052 7076
rect 75819 7027 75861 7036
rect 75436 6952 75572 6992
rect 74859 6572 74901 6581
rect 74859 6532 74860 6572
rect 74900 6532 74901 6572
rect 74859 6523 74901 6532
rect 74763 6320 74805 6329
rect 74763 6280 74764 6320
rect 74804 6280 74805 6320
rect 74763 6271 74805 6280
rect 74380 6236 74420 6245
rect 74380 5657 74420 6196
rect 74764 6186 74804 6271
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 74379 5648 74421 5657
rect 74379 5608 74380 5648
rect 74420 5608 74421 5648
rect 74379 5599 74421 5608
rect 74764 5648 74804 5657
rect 74475 4808 74517 4817
rect 74475 4768 74476 4808
rect 74516 4768 74517 4808
rect 74475 4759 74517 4768
rect 74476 4674 74516 4759
rect 73707 4304 73749 4313
rect 73707 4264 73708 4304
rect 73748 4264 73749 4304
rect 73707 4255 73749 4264
rect 74283 4304 74325 4313
rect 74283 4264 74284 4304
rect 74324 4264 74325 4304
rect 74283 4255 74325 4264
rect 73132 4136 73172 4145
rect 73132 3473 73172 4096
rect 73708 3557 73748 4255
rect 74284 4170 74324 4255
rect 74475 4220 74517 4229
rect 74475 4180 74476 4220
rect 74516 4180 74517 4220
rect 74475 4171 74517 4180
rect 74476 4136 74516 4171
rect 74764 4145 74804 5608
rect 75532 5396 75572 6952
rect 75819 6824 75861 6833
rect 75819 6784 75820 6824
rect 75860 6784 75861 6824
rect 75819 6775 75861 6784
rect 75628 6497 75668 6582
rect 75723 6572 75765 6581
rect 75723 6532 75724 6572
rect 75764 6532 75765 6572
rect 75723 6523 75765 6532
rect 75627 6488 75669 6497
rect 75627 6448 75628 6488
rect 75668 6448 75669 6488
rect 75627 6439 75669 6448
rect 75724 6488 75764 6523
rect 75724 6437 75764 6448
rect 75820 6488 75860 6775
rect 76012 6572 76052 7036
rect 76107 7036 76108 7076
rect 76148 7036 76149 7076
rect 76107 7027 76149 7036
rect 76300 6992 76340 7120
rect 76683 7160 76725 7169
rect 76683 7120 76684 7160
rect 76724 7120 76725 7160
rect 76683 7111 76725 7120
rect 76204 6952 76340 6992
rect 76204 6656 76244 6952
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 76204 6616 76340 6656
rect 76012 6532 76244 6572
rect 75820 6439 75860 6448
rect 75916 6488 75956 6497
rect 76204 6488 76244 6532
rect 76300 6497 76340 6616
rect 76491 6572 76533 6581
rect 76491 6532 76492 6572
rect 76532 6532 76533 6572
rect 76491 6523 76533 6532
rect 75956 6448 76148 6488
rect 75916 6439 75956 6448
rect 75627 6320 75669 6329
rect 75627 6280 75628 6320
rect 75668 6280 75669 6320
rect 75627 6271 75669 6280
rect 75628 5648 75668 6271
rect 76108 5648 76148 6448
rect 76204 6439 76244 6448
rect 76299 6488 76341 6497
rect 76299 6448 76300 6488
rect 76340 6448 76341 6488
rect 76299 6439 76341 6448
rect 76492 6488 76532 6523
rect 76492 6437 76532 6448
rect 76587 6488 76629 6497
rect 76587 6448 76588 6488
rect 76628 6448 76629 6488
rect 76587 6439 76629 6448
rect 76588 6354 76628 6439
rect 76204 5648 76244 5657
rect 76108 5608 76204 5648
rect 75628 5599 75668 5608
rect 76204 5599 76244 5608
rect 76395 5648 76437 5657
rect 76395 5608 76396 5648
rect 76436 5608 76437 5648
rect 76395 5599 76437 5608
rect 76492 5648 76532 5657
rect 76780 5648 76820 7792
rect 77164 7664 77204 7960
rect 77259 8000 77301 8009
rect 77259 7960 77260 8000
rect 77300 7960 77301 8000
rect 77259 7951 77301 7960
rect 77260 7866 77300 7951
rect 77356 7748 77396 9127
rect 77452 8672 77492 8681
rect 77452 7832 77492 8632
rect 78028 8009 78068 9220
rect 78316 8672 78356 10135
rect 78027 8000 78069 8009
rect 78027 7960 78028 8000
rect 78068 7960 78069 8000
rect 78027 7951 78069 7960
rect 77740 7832 77780 7841
rect 77452 7792 77740 7832
rect 77740 7783 77780 7792
rect 77356 7708 77492 7748
rect 77164 7624 77300 7664
rect 77163 7244 77205 7253
rect 77163 7204 77164 7244
rect 77204 7204 77205 7244
rect 77163 7195 77205 7204
rect 76972 7160 77012 7169
rect 76876 6320 76916 6329
rect 76972 6320 77012 7120
rect 77164 7160 77204 7195
rect 77260 7169 77300 7624
rect 77355 7328 77397 7337
rect 77355 7288 77356 7328
rect 77396 7288 77397 7328
rect 77355 7279 77397 7288
rect 77164 7109 77204 7120
rect 77259 7160 77301 7169
rect 77259 7120 77260 7160
rect 77300 7120 77301 7160
rect 77259 7111 77301 7120
rect 77068 7076 77108 7085
rect 77068 6656 77108 7036
rect 77068 6616 77300 6656
rect 76916 6280 77012 6320
rect 77068 6488 77108 6497
rect 76876 6271 76916 6280
rect 77068 5900 77108 6448
rect 77164 5900 77204 5909
rect 77068 5860 77164 5900
rect 77164 5851 77204 5860
rect 77260 5657 77300 6616
rect 77356 6488 77396 7279
rect 77452 7160 77492 7708
rect 77835 7328 77877 7337
rect 77835 7288 77836 7328
rect 77876 7288 77877 7328
rect 77835 7279 77877 7288
rect 77836 7194 77876 7279
rect 77452 7111 77492 7120
rect 77643 7160 77685 7169
rect 77643 7120 77644 7160
rect 77684 7120 77685 7160
rect 77643 7111 77685 7120
rect 77548 7076 77588 7085
rect 77452 6488 77492 6497
rect 77356 6448 77452 6488
rect 77452 6439 77492 6448
rect 77164 5648 77204 5657
rect 76780 5608 77164 5648
rect 76012 5564 76052 5573
rect 76012 5480 76052 5524
rect 76396 5514 76436 5599
rect 76492 5489 76532 5608
rect 77164 5599 77204 5608
rect 77259 5648 77301 5657
rect 77356 5648 77396 5657
rect 77259 5608 77260 5648
rect 77300 5608 77356 5648
rect 77259 5599 77301 5608
rect 77356 5599 77396 5608
rect 77452 5648 77492 5657
rect 77548 5648 77588 7036
rect 77644 6581 77684 7111
rect 77643 6572 77685 6581
rect 77643 6532 77644 6572
rect 77684 6532 77685 6572
rect 77643 6523 77685 6532
rect 78316 6488 78356 8632
rect 78316 6439 78356 6448
rect 77492 5608 77588 5648
rect 77452 5599 77492 5608
rect 77260 5514 77300 5599
rect 76300 5480 76340 5489
rect 76012 5440 76300 5480
rect 76300 5431 76340 5440
rect 76491 5480 76533 5489
rect 76491 5440 76492 5480
rect 76532 5440 76533 5480
rect 76491 5431 76533 5440
rect 75532 5356 76052 5396
rect 75916 4976 75956 4985
rect 74859 4808 74901 4817
rect 74859 4768 74860 4808
rect 74900 4768 74901 4808
rect 74859 4759 74901 4768
rect 74476 4085 74516 4096
rect 74571 4136 74613 4145
rect 74571 4096 74572 4136
rect 74612 4096 74613 4136
rect 74571 4087 74613 4096
rect 74763 4136 74805 4145
rect 74763 4096 74764 4136
rect 74804 4096 74805 4136
rect 74763 4087 74805 4096
rect 74860 4136 74900 4759
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 75819 4304 75861 4313
rect 75916 4304 75956 4936
rect 76012 4976 76052 5356
rect 76107 5312 76149 5321
rect 76107 5272 76108 5312
rect 76148 5272 76149 5312
rect 76107 5263 76149 5272
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 76108 5144 76148 5263
rect 76108 5095 76148 5104
rect 76012 4304 76052 4936
rect 76204 4976 76244 4985
rect 76396 4976 76436 4985
rect 76204 4397 76244 4936
rect 76300 4936 76396 4976
rect 76203 4388 76245 4397
rect 76203 4348 76204 4388
rect 76244 4348 76245 4388
rect 76203 4339 76245 4348
rect 75819 4264 75820 4304
rect 75860 4264 75956 4304
rect 76009 4264 76052 4304
rect 75819 4255 75861 4264
rect 74860 4087 74900 4096
rect 75723 4136 75765 4145
rect 75723 4096 75724 4136
rect 75764 4096 75765 4136
rect 75723 4087 75765 4096
rect 73707 3548 73749 3557
rect 73707 3508 73708 3548
rect 73748 3508 73749 3548
rect 73707 3499 73749 3508
rect 74572 3473 74612 4087
rect 75724 4002 75764 4087
rect 75820 3557 75860 4255
rect 76009 4220 76049 4264
rect 76300 4220 76340 4936
rect 76396 4927 76436 4936
rect 76587 4976 76629 4985
rect 76587 4936 76588 4976
rect 76628 4936 76629 4976
rect 76587 4927 76629 4936
rect 76684 4976 76724 4985
rect 77164 4976 77204 4985
rect 76588 4842 76628 4927
rect 76396 4724 76436 4733
rect 76396 4229 76436 4684
rect 76684 4388 76724 4936
rect 76492 4348 76724 4388
rect 76972 4936 77164 4976
rect 76009 4180 76053 4220
rect 76013 4136 76053 4180
rect 76012 4096 76053 4136
rect 76108 4180 76340 4220
rect 76395 4220 76437 4229
rect 76395 4180 76396 4220
rect 76436 4180 76437 4220
rect 76012 3641 76052 4096
rect 76108 3884 76148 4180
rect 76395 4171 76437 4180
rect 76492 4052 76532 4348
rect 76875 4304 76917 4313
rect 76875 4264 76876 4304
rect 76916 4264 76917 4304
rect 76875 4255 76917 4264
rect 76876 4170 76916 4255
rect 76779 4136 76821 4145
rect 76779 4096 76780 4136
rect 76820 4096 76821 4136
rect 76779 4087 76821 4096
rect 76107 3844 76148 3884
rect 76204 4012 76532 4052
rect 76107 3716 76147 3844
rect 76107 3676 76148 3716
rect 76011 3632 76053 3641
rect 76011 3592 76012 3632
rect 76052 3592 76053 3632
rect 76011 3583 76053 3592
rect 76108 3632 76148 3676
rect 76108 3583 76148 3592
rect 75819 3548 75861 3557
rect 75819 3508 75820 3548
rect 75860 3508 75861 3548
rect 75819 3499 75861 3508
rect 72652 2827 72692 2836
rect 72075 2708 72117 2717
rect 72075 2668 72076 2708
rect 72116 2668 72117 2708
rect 72075 2659 72117 2668
rect 72076 2465 72116 2659
rect 72171 2624 72213 2633
rect 72171 2584 72172 2624
rect 72212 2584 72213 2624
rect 72171 2575 72213 2584
rect 72172 2490 72212 2575
rect 72075 2456 72117 2465
rect 72652 2456 72692 2465
rect 72075 2416 72076 2456
rect 72116 2416 72117 2456
rect 72075 2407 72117 2416
rect 72556 2416 72652 2456
rect 71924 1324 72020 1364
rect 71884 1315 71924 1324
rect 69388 1231 69428 1240
rect 68948 1072 69044 1112
rect 70731 1112 70773 1121
rect 70731 1072 70732 1112
rect 70772 1072 70773 1112
rect 68908 1063 68948 1072
rect 70731 1063 70773 1072
rect 71211 1112 71253 1121
rect 71211 1072 71212 1112
rect 71252 1072 71253 1112
rect 71211 1063 71253 1072
rect 72556 1112 72596 2416
rect 72652 2407 72692 2416
rect 72652 1952 72692 1961
rect 72748 1952 72788 3415
rect 72844 3221 72884 3424
rect 73036 3464 73076 3473
rect 72843 3212 72885 3221
rect 72843 3172 72844 3212
rect 72884 3172 72885 3212
rect 72843 3163 72885 3172
rect 72940 3212 72980 3221
rect 72940 2885 72980 3172
rect 73036 2900 73076 3424
rect 73131 3464 73173 3473
rect 73131 3424 73132 3464
rect 73172 3424 73173 3464
rect 73131 3415 73173 3424
rect 74571 3464 74613 3473
rect 74571 3424 74572 3464
rect 74612 3424 74613 3464
rect 74571 3415 74613 3424
rect 75820 3464 75860 3499
rect 73995 3296 74037 3305
rect 73995 3256 73996 3296
rect 74036 3256 74037 3296
rect 73995 3247 74037 3256
rect 72939 2876 72981 2885
rect 72939 2836 72940 2876
rect 72980 2836 72981 2876
rect 73036 2876 73364 2900
rect 73036 2860 73324 2876
rect 72939 2827 72981 2836
rect 73324 2827 73364 2836
rect 72940 2717 72980 2827
rect 73611 2792 73653 2801
rect 73611 2752 73612 2792
rect 73652 2752 73653 2792
rect 73611 2743 73653 2752
rect 73899 2792 73941 2801
rect 73899 2752 73900 2792
rect 73940 2752 73941 2792
rect 73899 2743 73941 2752
rect 72939 2708 72981 2717
rect 72939 2668 72940 2708
rect 72980 2668 72981 2708
rect 72939 2659 72981 2668
rect 73612 2624 73652 2743
rect 73612 2120 73652 2584
rect 73707 2624 73749 2633
rect 73707 2584 73708 2624
rect 73748 2584 73749 2624
rect 73707 2575 73749 2584
rect 73708 2490 73748 2575
rect 73804 2120 73844 2129
rect 73612 2080 73804 2120
rect 73804 1961 73844 2080
rect 72692 1912 72788 1952
rect 73803 1952 73845 1961
rect 73803 1912 73804 1952
rect 73844 1912 73845 1952
rect 72652 1903 72692 1912
rect 73803 1903 73845 1912
rect 72556 1063 72596 1072
rect 73227 1112 73269 1121
rect 73227 1072 73228 1112
rect 73268 1072 73269 1112
rect 73227 1063 73269 1072
rect 73612 1112 73652 1121
rect 73900 1112 73940 2743
rect 73996 2624 74036 3247
rect 74187 2708 74229 2717
rect 74187 2668 74188 2708
rect 74228 2668 74229 2708
rect 74187 2659 74229 2668
rect 74475 2708 74517 2717
rect 74475 2668 74476 2708
rect 74516 2668 74517 2708
rect 74475 2659 74517 2668
rect 73996 2549 74036 2584
rect 73995 2540 74037 2549
rect 73995 2500 73996 2540
rect 74036 2500 74037 2540
rect 73995 2491 74037 2500
rect 73995 2204 74037 2213
rect 73995 2164 73996 2204
rect 74036 2164 74037 2204
rect 73995 2155 74037 2164
rect 73996 1952 74036 2155
rect 73996 1877 74036 1912
rect 74188 1952 74228 2659
rect 74283 2624 74325 2633
rect 74283 2584 74284 2624
rect 74324 2584 74325 2624
rect 74283 2575 74325 2584
rect 74476 2624 74516 2659
rect 74284 2490 74324 2575
rect 74380 2540 74420 2549
rect 74188 1903 74228 1912
rect 74284 1952 74324 1961
rect 74380 1952 74420 2500
rect 74476 2297 74516 2584
rect 74475 2288 74517 2297
rect 74475 2248 74476 2288
rect 74516 2248 74517 2288
rect 74475 2239 74517 2248
rect 74572 2120 74612 3415
rect 75820 3414 75860 3424
rect 75916 3464 75956 3473
rect 74859 3380 74901 3389
rect 74859 3340 74860 3380
rect 74900 3340 74901 3380
rect 74859 3331 74901 3340
rect 74860 2969 74900 3331
rect 75916 3212 75956 3424
rect 75820 3172 75956 3212
rect 76012 3464 76052 3473
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 74859 2960 74901 2969
rect 74859 2920 74860 2960
rect 74900 2920 74901 2960
rect 74859 2911 74901 2920
rect 74667 2792 74709 2801
rect 74667 2752 74668 2792
rect 74708 2752 74709 2792
rect 74667 2743 74709 2752
rect 74668 2658 74708 2743
rect 74763 2624 74805 2633
rect 74763 2584 74764 2624
rect 74804 2584 74805 2624
rect 74763 2575 74805 2584
rect 74667 2288 74709 2297
rect 74667 2248 74668 2288
rect 74708 2248 74709 2288
rect 74667 2239 74709 2248
rect 74324 1912 74420 1952
rect 74476 2080 74612 2120
rect 74284 1903 74324 1912
rect 73995 1868 74037 1877
rect 73995 1828 73996 1868
rect 74036 1828 74037 1868
rect 73995 1819 74037 1828
rect 73996 1700 74036 1709
rect 73996 1121 74036 1660
rect 73652 1072 73940 1112
rect 73995 1112 74037 1121
rect 73995 1072 73996 1112
rect 74036 1072 74037 1112
rect 73612 1063 73652 1072
rect 73995 1063 74037 1072
rect 74476 1112 74516 2080
rect 74571 1952 74613 1961
rect 74571 1912 74572 1952
rect 74612 1912 74613 1952
rect 74571 1903 74613 1912
rect 74668 1952 74708 2239
rect 74668 1903 74708 1912
rect 74572 1818 74612 1903
rect 74764 1625 74804 2575
rect 74860 1952 74900 2911
rect 75820 2465 75860 3172
rect 76012 3137 76052 3424
rect 76107 3464 76149 3473
rect 76107 3424 76108 3464
rect 76148 3424 76149 3464
rect 76107 3415 76149 3424
rect 76011 3128 76053 3137
rect 75916 3088 76012 3128
rect 76052 3088 76053 3128
rect 75819 2456 75861 2465
rect 75819 2416 75820 2456
rect 75860 2416 75861 2456
rect 75819 2407 75861 2416
rect 75436 2080 75860 2120
rect 74860 1903 74900 1912
rect 75148 1952 75188 1961
rect 74860 1784 74900 1793
rect 75148 1784 75188 1912
rect 75243 1952 75285 1961
rect 75243 1912 75244 1952
rect 75284 1912 75285 1952
rect 75243 1903 75285 1912
rect 75436 1952 75476 2080
rect 75436 1903 75476 1912
rect 75628 1952 75668 1961
rect 75244 1818 75284 1903
rect 74900 1744 75188 1784
rect 75436 1784 75476 1793
rect 75628 1784 75668 1912
rect 75476 1744 75668 1784
rect 74860 1735 74900 1744
rect 75436 1735 75476 1744
rect 74763 1616 74805 1625
rect 74763 1576 74764 1616
rect 74804 1576 74805 1616
rect 74763 1567 74805 1576
rect 75627 1616 75669 1625
rect 75627 1576 75628 1616
rect 75668 1576 75669 1616
rect 75627 1567 75669 1576
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 75628 1364 75668 1567
rect 75628 1315 75668 1324
rect 74476 1063 74516 1072
rect 70732 978 70772 1063
rect 71212 978 71252 1063
rect 73228 978 73268 1063
rect 68524 904 68756 944
rect 75820 944 75860 2080
rect 75916 1112 75956 3088
rect 76011 3079 76053 3088
rect 76108 2969 76148 3415
rect 76107 2960 76149 2969
rect 76107 2920 76108 2960
rect 76148 2920 76149 2960
rect 76107 2911 76149 2920
rect 76012 2792 76052 2801
rect 76012 1952 76052 2752
rect 76108 2624 76148 2911
rect 76204 2876 76244 4012
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 76780 3716 76820 4087
rect 76780 3676 76916 3716
rect 76299 3632 76341 3641
rect 76299 3592 76300 3632
rect 76340 3592 76341 3632
rect 76299 3583 76341 3592
rect 76204 2827 76244 2836
rect 76300 2708 76340 3583
rect 76779 3548 76821 3557
rect 76779 3508 76780 3548
rect 76820 3508 76821 3548
rect 76779 3499 76821 3508
rect 76396 3464 76436 3473
rect 76396 3305 76436 3424
rect 76683 3464 76725 3473
rect 76683 3424 76684 3464
rect 76724 3424 76725 3464
rect 76683 3415 76725 3424
rect 76684 3330 76724 3415
rect 76780 3414 76820 3499
rect 76395 3296 76437 3305
rect 76395 3256 76396 3296
rect 76436 3256 76437 3296
rect 76395 3247 76437 3256
rect 76779 3296 76821 3305
rect 76779 3256 76780 3296
rect 76820 3256 76821 3296
rect 76779 3247 76821 3256
rect 76395 2708 76437 2717
rect 76300 2668 76396 2708
rect 76436 2668 76437 2708
rect 76395 2659 76437 2668
rect 76204 2624 76244 2633
rect 76108 2584 76204 2624
rect 76204 2575 76244 2584
rect 76396 2624 76436 2659
rect 76396 2573 76436 2584
rect 76492 2624 76532 2633
rect 76780 2624 76820 3247
rect 76876 2969 76916 3676
rect 76875 2960 76917 2969
rect 76875 2920 76876 2960
rect 76916 2920 76917 2960
rect 76875 2911 76917 2920
rect 76532 2584 76628 2624
rect 76492 2575 76532 2584
rect 76107 2456 76149 2465
rect 76107 2416 76108 2456
rect 76148 2416 76149 2456
rect 76588 2456 76628 2584
rect 76780 2575 76820 2584
rect 76779 2456 76821 2465
rect 76588 2416 76780 2456
rect 76820 2416 76821 2456
rect 76107 2407 76149 2416
rect 76779 2407 76821 2416
rect 76012 1903 76052 1912
rect 76012 1112 76052 1121
rect 75916 1072 76012 1112
rect 76012 1063 76052 1072
rect 76108 1112 76148 2407
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 76780 1121 76820 2407
rect 76876 1952 76916 2911
rect 76972 2213 77012 4936
rect 77164 4927 77204 4936
rect 77355 4976 77397 4985
rect 77355 4936 77356 4976
rect 77396 4936 77397 4976
rect 77355 4927 77397 4936
rect 77452 4976 77492 4985
rect 77492 4936 77780 4976
rect 77452 4927 77492 4936
rect 77164 4724 77204 4733
rect 77068 4684 77164 4724
rect 77068 4136 77108 4684
rect 77164 4675 77204 4684
rect 77068 4087 77108 4096
rect 77356 3548 77396 4927
rect 77451 4808 77493 4817
rect 77451 4768 77452 4808
rect 77492 4768 77493 4808
rect 77451 4759 77493 4768
rect 77452 4136 77492 4759
rect 77452 4087 77492 4096
rect 77356 3499 77396 3508
rect 77740 3548 77780 4936
rect 77835 4808 77877 4817
rect 77835 4768 77836 4808
rect 77876 4768 77877 4808
rect 77835 4759 77877 4768
rect 77836 4674 77876 4759
rect 78412 4313 78452 15763
rect 78603 14972 78645 14981
rect 78603 14932 78604 14972
rect 78644 14932 78645 14972
rect 78603 14923 78645 14932
rect 78604 14838 78644 14923
rect 78603 14552 78645 14561
rect 78603 14512 78604 14552
rect 78644 14512 78645 14552
rect 78603 14503 78645 14512
rect 78604 14418 78644 14503
rect 78700 14225 78740 16192
rect 78891 16192 78892 16232
rect 78932 16192 78933 16232
rect 78891 16183 78933 16192
rect 79180 16232 79220 17032
rect 79276 16484 79316 17116
rect 79371 17116 79372 17156
rect 79412 17116 79413 17156
rect 79371 17107 79413 17116
rect 79276 16435 79316 16444
rect 78892 16098 78932 16183
rect 79180 14981 79220 16192
rect 79372 15560 79412 17107
rect 79545 17072 79585 17472
rect 79655 17165 79695 17472
rect 79654 17156 79696 17165
rect 79654 17116 79655 17156
rect 79695 17116 79696 17156
rect 79654 17107 79696 17116
rect 79468 17032 79585 17072
rect 79468 15728 79508 17032
rect 79468 15679 79508 15688
rect 79372 15511 79412 15520
rect 79179 14972 79221 14981
rect 79179 14932 79180 14972
rect 79220 14932 79221 14972
rect 79179 14923 79221 14932
rect 78699 14216 78741 14225
rect 78699 14176 78700 14216
rect 78740 14176 78741 14216
rect 78699 14167 78741 14176
rect 79371 14216 79413 14225
rect 79371 14176 79372 14216
rect 79412 14176 79413 14216
rect 79371 14167 79413 14176
rect 79372 14082 79412 14167
rect 79275 12284 79317 12293
rect 79275 12244 79276 12284
rect 79316 12244 79317 12284
rect 79275 12235 79317 12244
rect 79276 12150 79316 12235
rect 79467 10268 79509 10277
rect 79467 10228 79468 10268
rect 79508 10228 79509 10268
rect 79467 10219 79509 10228
rect 79468 10134 79508 10219
rect 79467 9680 79509 9689
rect 79467 9640 79468 9680
rect 79508 9640 79509 9680
rect 79467 9631 79509 9640
rect 79468 8924 79508 9631
rect 79468 8875 79508 8884
rect 79468 6656 79508 6667
rect 79468 6581 79508 6616
rect 79467 6572 79509 6581
rect 79467 6532 79468 6572
rect 79508 6532 79509 6572
rect 79467 6523 79509 6532
rect 77835 4304 77877 4313
rect 77835 4264 77836 4304
rect 77876 4264 77877 4304
rect 77835 4255 77877 4264
rect 78411 4304 78453 4313
rect 78411 4264 78412 4304
rect 78452 4264 78453 4304
rect 78411 4255 78453 4264
rect 79467 4304 79509 4313
rect 79467 4264 79468 4304
rect 79508 4264 79509 4304
rect 79467 4255 79509 4264
rect 77740 3499 77780 3508
rect 77836 3473 77876 4255
rect 79468 4170 79508 4255
rect 78316 4136 78356 4145
rect 77260 3464 77300 3473
rect 77068 3296 77108 3305
rect 77260 3296 77300 3424
rect 77108 3256 77300 3296
rect 77452 3464 77492 3473
rect 77068 3247 77108 3256
rect 77452 3221 77492 3424
rect 77644 3464 77684 3473
rect 77451 3212 77493 3221
rect 77451 3172 77452 3212
rect 77492 3172 77493 3212
rect 77451 3163 77493 3172
rect 77644 2900 77684 3424
rect 77835 3464 77877 3473
rect 77835 3424 77836 3464
rect 77876 3424 77877 3464
rect 77835 3415 77877 3424
rect 77836 3330 77876 3415
rect 77835 3212 77877 3221
rect 77835 3172 77836 3212
rect 77876 3172 77877 3212
rect 77835 3163 77877 3172
rect 77356 2860 77684 2900
rect 77356 2717 77396 2860
rect 77452 2792 77492 2801
rect 77492 2752 77684 2792
rect 77452 2743 77492 2752
rect 77355 2708 77397 2717
rect 77355 2668 77356 2708
rect 77396 2668 77397 2708
rect 77355 2659 77397 2668
rect 77067 2624 77109 2633
rect 77067 2584 77068 2624
rect 77108 2584 77109 2624
rect 77067 2575 77109 2584
rect 76971 2204 77013 2213
rect 76971 2164 76972 2204
rect 77012 2164 77013 2204
rect 76971 2155 77013 2164
rect 76876 1903 76916 1912
rect 77068 1364 77108 2575
rect 77164 2540 77204 2551
rect 77164 2465 77204 2500
rect 77356 2465 77396 2659
rect 77644 2624 77684 2752
rect 77644 2575 77684 2584
rect 77836 2624 77876 3163
rect 78316 2969 78356 4096
rect 78123 2960 78165 2969
rect 78123 2920 78124 2960
rect 78164 2920 78165 2960
rect 78123 2911 78165 2920
rect 78315 2960 78357 2969
rect 78315 2920 78316 2960
rect 78356 2920 78357 2960
rect 78315 2911 78357 2920
rect 77836 2575 77876 2584
rect 77740 2540 77780 2549
rect 77163 2456 77205 2465
rect 77163 2416 77164 2456
rect 77204 2416 77205 2456
rect 77163 2407 77205 2416
rect 77355 2456 77397 2465
rect 77355 2416 77356 2456
rect 77396 2416 77397 2456
rect 77355 2407 77397 2416
rect 77740 1961 77780 2500
rect 77739 1952 77781 1961
rect 77739 1912 77740 1952
rect 77780 1912 77781 1952
rect 77739 1903 77781 1912
rect 77068 1315 77108 1324
rect 78028 1700 78068 1709
rect 78028 1121 78068 1660
rect 76108 1063 76148 1072
rect 76203 1112 76245 1121
rect 76203 1072 76204 1112
rect 76244 1072 76245 1112
rect 76203 1063 76245 1072
rect 76779 1112 76821 1121
rect 76779 1072 76780 1112
rect 76820 1072 76821 1112
rect 76779 1063 76821 1072
rect 78027 1112 78069 1121
rect 78027 1072 78028 1112
rect 78068 1072 78069 1112
rect 78124 1112 78164 2911
rect 78220 2792 78260 2801
rect 78260 2752 78356 2792
rect 78220 2743 78260 2752
rect 78219 2204 78261 2213
rect 78219 2164 78220 2204
rect 78260 2164 78261 2204
rect 78219 2155 78261 2164
rect 78220 1952 78260 2155
rect 78220 1903 78260 1912
rect 78220 1700 78260 1709
rect 78220 1289 78260 1660
rect 78219 1280 78261 1289
rect 78219 1240 78220 1280
rect 78260 1240 78261 1280
rect 78219 1231 78261 1240
rect 78220 1112 78260 1121
rect 78124 1072 78220 1112
rect 78316 1112 78356 2752
rect 78891 2624 78933 2633
rect 78891 2584 78892 2624
rect 78932 2584 78933 2624
rect 78891 2575 78933 2584
rect 78699 2456 78741 2465
rect 78699 2416 78700 2456
rect 78740 2416 78741 2456
rect 78699 2407 78741 2416
rect 78411 1952 78453 1961
rect 78411 1912 78412 1952
rect 78452 1912 78453 1952
rect 78411 1903 78453 1912
rect 78508 1952 78548 1961
rect 78412 1818 78452 1903
rect 78508 1784 78548 1912
rect 78700 1952 78740 2407
rect 78700 1903 78740 1912
rect 78892 1952 78932 2575
rect 78892 1903 78932 1912
rect 78796 1784 78836 1793
rect 78508 1744 78796 1784
rect 78796 1735 78836 1744
rect 79467 1280 79509 1289
rect 79467 1240 79468 1280
rect 79508 1240 79509 1280
rect 79467 1231 79509 1240
rect 79084 1112 79124 1121
rect 78316 1072 79084 1112
rect 78027 1063 78069 1072
rect 78220 1063 78260 1072
rect 79084 1063 79124 1072
rect 79468 1112 79508 1231
rect 79468 1063 79508 1072
rect 76204 978 76244 1063
rect 75916 944 75956 953
rect 75820 904 75916 944
rect 64203 895 64245 904
rect 75916 895 75956 904
rect 57004 820 57332 860
rect 60364 810 60404 895
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 652 37528 692 37568
rect 55948 37948 55988 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 844 25936 884 25976
rect 652 25768 692 25808
rect 844 25096 884 25136
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 844 23836 884 23876
rect 844 23584 884 23624
rect 652 23248 692 23288
rect 556 22408 596 22448
rect 652 21568 692 21608
rect 844 21568 884 21608
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 54412 36772 54452 36812
rect 38668 36688 38708 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 3820 30556 3860 30596
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 38476 28540 38516 28580
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 37804 27700 37844 27740
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 2764 25096 2804 25136
rect 1804 24004 1844 24044
rect 2188 24004 2228 24044
rect 1996 23836 2036 23876
rect 1420 23584 1460 23624
rect 1516 23164 1556 23204
rect 1420 23080 1460 23120
rect 1900 23080 1940 23120
rect 2092 23080 2132 23120
rect 940 21400 980 21440
rect 1708 21316 1748 21356
rect 652 20728 692 20768
rect 1900 22324 1940 22364
rect 2668 21316 2708 21356
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 1708 17788 1748 17828
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 844 15436 884 15476
rect 652 14848 692 14888
rect 1036 14932 1076 14972
rect 1708 17200 1748 17240
rect 1036 14008 1076 14048
rect 1324 13924 1364 13964
rect 748 13756 788 13796
rect 652 13168 692 13208
rect 652 12328 692 12368
rect 652 11488 692 11528
rect 652 10732 692 10772
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 1516 14680 1556 14720
rect 2476 17200 2516 17240
rect 2668 16948 2708 16988
rect 2380 16360 2420 16400
rect 2188 15940 2228 15980
rect 2188 15688 2228 15728
rect 1996 14932 2036 14972
rect 1804 14848 1844 14888
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3628 23080 3668 23120
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3244 22324 3284 22364
rect 3244 21736 3284 21776
rect 3052 21568 3092 21608
rect 3148 21400 3188 21440
rect 3244 21316 3284 21356
rect 3532 21316 3572 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 33484 26188 33524 26228
rect 34252 26188 34292 26228
rect 32716 26104 32756 26144
rect 31948 25936 31988 25976
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 29836 24676 29876 24716
rect 33964 26104 34004 26144
rect 33484 25936 33524 25976
rect 33148 25852 33188 25892
rect 31084 24508 31124 24548
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 28204 23164 28244 23204
rect 3820 23080 3860 23120
rect 2860 21064 2900 21104
rect 3628 21064 3668 21104
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 29548 23836 29588 23876
rect 22060 22996 22100 23036
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 5548 21400 5588 21440
rect 4780 21316 4820 21356
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 5932 21484 5972 21524
rect 5740 21316 5780 21356
rect 6124 21316 6164 21356
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 6124 20728 6164 20768
rect 4780 18376 4820 18416
rect 3916 18124 3956 18164
rect 3820 18040 3860 18080
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 2572 16108 2612 16148
rect 2956 16108 2996 16148
rect 2668 15940 2708 15980
rect 1612 14260 1652 14300
rect 2188 14260 2228 14300
rect 1516 13756 1556 13796
rect 1420 13000 1460 13040
rect 1324 12412 1364 12452
rect 1324 12160 1364 12200
rect 1708 13168 1748 13208
rect 2380 14260 2420 14300
rect 2284 14176 2324 14216
rect 2380 13504 2420 13544
rect 2092 12580 2132 12620
rect 3628 16024 3668 16064
rect 3436 15688 3476 15728
rect 2956 15268 2996 15308
rect 3436 15268 3476 15308
rect 2860 15100 2900 15140
rect 2764 14848 2804 14888
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 2956 14680 2996 14720
rect 2956 14428 2996 14468
rect 2860 14176 2900 14216
rect 2764 13504 2804 13544
rect 2476 13336 2516 13376
rect 2764 13336 2804 13376
rect 1612 12328 1652 12368
rect 1516 12244 1556 12284
rect 1900 12244 1940 12284
rect 2572 12664 2612 12704
rect 2284 12328 2324 12368
rect 2476 12328 2516 12368
rect 2188 12244 2228 12284
rect 1708 12160 1748 12200
rect 1996 12160 2036 12200
rect 1420 11740 1460 11780
rect 940 10312 980 10352
rect 844 9640 884 9680
rect 844 9388 884 9428
rect 1324 10396 1364 10436
rect 2092 11824 2132 11864
rect 1996 11656 2036 11696
rect 1516 10312 1556 10352
rect 1612 10228 1652 10268
rect 2668 11656 2708 11696
rect 2188 10312 2228 10352
rect 3052 14008 3092 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 3340 13336 3380 13376
rect 3340 13084 3380 13124
rect 3628 13000 3668 13040
rect 2956 12664 2996 12704
rect 2860 12328 2900 12368
rect 2476 10312 2516 10352
rect 2380 10144 2420 10184
rect 1516 9640 1556 9680
rect 1420 9388 1460 9428
rect 652 8128 692 8168
rect 652 7288 692 7328
rect 1708 8632 1748 8672
rect 1228 8548 1268 8588
rect 1132 8128 1172 8168
rect 1996 9472 2036 9512
rect 1996 8716 2036 8756
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 1036 7540 1076 7580
rect 1228 5524 1268 5564
rect 1804 7960 1844 8000
rect 1804 7540 1844 7580
rect 1516 6616 1556 6656
rect 1516 5692 1556 5732
rect 1420 5440 1460 5480
rect 1708 5440 1748 5480
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3436 11908 3476 11948
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4204 16444 4244 16484
rect 4012 16360 4052 16400
rect 3916 14260 3956 14300
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 5548 19972 5588 20012
rect 9004 19972 9044 20012
rect 6604 19384 6644 19424
rect 7948 19384 7988 19424
rect 8812 19384 8852 19424
rect 5932 17620 5972 17660
rect 5452 16948 5492 16988
rect 4876 16444 4916 16484
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4300 15688 4340 15728
rect 4204 15520 4244 15560
rect 4780 15520 4820 15560
rect 4684 15436 4724 15476
rect 4492 15352 4532 15392
rect 5836 16192 5876 16232
rect 8524 19300 8564 19340
rect 9004 19300 9044 19340
rect 8332 18880 8372 18920
rect 8620 19216 8660 19256
rect 9100 19216 9140 19256
rect 8812 18880 8852 18920
rect 8524 18796 8564 18836
rect 8908 18796 8948 18836
rect 8044 18544 8084 18584
rect 8524 18544 8564 18584
rect 7948 17788 7988 17828
rect 8620 18124 8660 18164
rect 8620 17956 8660 17996
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 21964 19552 22004 19592
rect 11692 19468 11732 19508
rect 9292 19384 9332 19424
rect 21580 19300 21620 19340
rect 9484 19216 9524 19256
rect 9196 18628 9236 18668
rect 8908 17956 8948 17996
rect 8044 17620 8084 17660
rect 7660 16360 7700 16400
rect 6316 16192 6356 16232
rect 7084 16192 7124 16232
rect 4780 14596 4820 14636
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4300 14092 4340 14132
rect 3340 11824 3380 11864
rect 3532 11824 3572 11864
rect 3436 11404 3476 11444
rect 2668 10312 2708 10352
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3436 10396 3476 10436
rect 2476 8464 2516 8504
rect 2380 8128 2420 8168
rect 2860 10060 2900 10100
rect 2860 9640 2900 9680
rect 3340 10228 3380 10268
rect 3148 10060 3188 10100
rect 2956 9472 2996 9512
rect 3244 9472 3284 9512
rect 3148 9388 3188 9428
rect 4396 14008 4436 14048
rect 4300 13924 4340 13964
rect 4684 13756 4724 13796
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 4588 12664 4628 12704
rect 4492 12496 4532 12536
rect 3724 11656 3764 11696
rect 3628 11572 3668 11612
rect 3628 11404 3668 11444
rect 3532 9640 3572 9680
rect 3916 11824 3956 11864
rect 3916 11656 3956 11696
rect 3820 11068 3860 11108
rect 3628 9556 3668 9596
rect 5260 14680 5300 14720
rect 5164 14596 5204 14636
rect 4876 14428 4916 14468
rect 5260 14092 5300 14132
rect 4876 13252 4916 13292
rect 5164 13168 5204 13208
rect 5068 12664 5108 12704
rect 4204 11488 4244 11528
rect 4684 11488 4724 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 5068 11572 5108 11612
rect 4588 11152 4628 11192
rect 4300 11068 4340 11108
rect 4204 10144 4244 10184
rect 4876 10984 4916 11024
rect 5068 10312 5108 10352
rect 4876 10228 4916 10268
rect 4588 9976 4628 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4492 9556 4532 9596
rect 4780 9556 4820 9596
rect 3436 9220 3476 9260
rect 2764 8800 2804 8840
rect 2572 7792 2612 7832
rect 3628 9220 3668 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3436 8800 3476 8840
rect 2764 7792 2804 7832
rect 2284 7036 2324 7076
rect 2188 6616 2228 6656
rect 3052 7960 3092 8000
rect 3532 8716 3572 8756
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2380 6280 2420 6320
rect 2572 6280 2612 6320
rect 2188 5524 2228 5564
rect 2284 5104 2324 5144
rect 2956 7120 2996 7160
rect 3820 8464 3860 8504
rect 3820 7960 3860 8000
rect 3724 7708 3764 7748
rect 4300 9472 4340 9512
rect 4492 9388 4532 9428
rect 4876 9472 4916 9512
rect 4588 9304 4628 9344
rect 4780 8800 4820 8840
rect 4492 8632 4532 8672
rect 5452 13336 5492 13376
rect 5356 13084 5396 13124
rect 5356 12328 5396 12368
rect 5260 10312 5300 10352
rect 4972 8800 5012 8840
rect 4972 8632 5012 8672
rect 4396 8464 4436 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4588 7960 4628 8000
rect 3628 6532 3668 6572
rect 3916 6532 3956 6572
rect 3532 6448 3572 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 2956 5692 2996 5732
rect 1036 3928 1076 3968
rect 1324 3508 1364 3548
rect 1132 3340 1172 3380
rect 3628 5692 3668 5732
rect 2764 5020 2804 5060
rect 1900 3256 1940 3296
rect 652 3088 692 3128
rect 1612 3172 1652 3212
rect 1708 2668 1748 2708
rect 2668 4012 2708 4052
rect 2572 3928 2612 3968
rect 3436 5272 3476 5312
rect 3532 5188 3572 5228
rect 3436 4936 3476 4976
rect 5164 7708 5204 7748
rect 4972 7120 5012 7160
rect 4300 7036 4340 7076
rect 4780 7036 4820 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 4204 6532 4244 6572
rect 4492 6448 4532 6488
rect 4204 6028 4244 6068
rect 4972 6028 5012 6068
rect 4108 5692 4148 5732
rect 4012 5272 4052 5312
rect 5068 5860 5108 5900
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3916 5104 3956 5144
rect 4300 5020 4340 5060
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 3052 4096 3092 4136
rect 2956 3508 2996 3548
rect 3820 4264 3860 4304
rect 3724 4012 3764 4052
rect 3916 4012 3956 4052
rect 3532 3928 3572 3968
rect 2476 3340 2516 3380
rect 2380 2584 2420 2624
rect 2668 3256 2708 3296
rect 2572 3172 2612 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 4684 4936 4724 4976
rect 4012 3928 4052 3968
rect 4396 4264 4436 4304
rect 4492 4180 4532 4220
rect 4588 3928 4628 3968
rect 5740 5608 5780 5648
rect 5740 5020 5780 5060
rect 6796 16024 6836 16064
rect 6988 16024 7028 16064
rect 6796 15856 6836 15896
rect 6220 13336 6260 13376
rect 6604 13756 6644 13796
rect 6700 13252 6740 13292
rect 8812 17200 8852 17240
rect 8716 15856 8756 15896
rect 6988 15436 7028 15476
rect 9580 18544 9620 18584
rect 10540 19216 10580 19256
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 11692 18544 11732 18584
rect 21484 18208 21524 18248
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 9580 17788 9620 17828
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 9388 16444 9428 16484
rect 21772 19048 21812 19088
rect 21868 18208 21908 18248
rect 21676 17704 21716 17744
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 27532 22156 27572 22196
rect 28012 22156 28052 22196
rect 22252 21652 22292 21692
rect 22156 19468 22196 19508
rect 25900 21484 25940 21524
rect 26860 21484 26900 21524
rect 22348 21316 22388 21356
rect 26476 21400 26516 21440
rect 27436 21316 27476 21356
rect 26860 21232 26900 21272
rect 25900 21064 25940 21104
rect 26668 20980 26708 21020
rect 24076 20224 24116 20264
rect 22540 19804 22580 19844
rect 22828 19804 22868 19844
rect 22060 18628 22100 18668
rect 22540 18880 22580 18920
rect 22540 18544 22580 18584
rect 22444 18460 22484 18500
rect 22252 18292 22292 18332
rect 22444 18292 22484 18332
rect 22444 17956 22484 17996
rect 22924 19048 22964 19088
rect 22828 18880 22868 18920
rect 22924 18712 22964 18752
rect 25804 20056 25844 20096
rect 25612 19972 25652 20012
rect 26284 19972 26324 20012
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 26956 20224 26996 20264
rect 27244 20224 27284 20264
rect 26764 19972 26804 20012
rect 23116 18628 23156 18668
rect 23020 18544 23060 18584
rect 22828 18460 22868 18500
rect 22732 17956 22772 17996
rect 22636 17872 22676 17912
rect 23020 18124 23060 18164
rect 22636 17704 22676 17744
rect 22828 17704 22868 17744
rect 22732 17620 22772 17660
rect 22540 17368 22580 17408
rect 22732 17368 22772 17408
rect 23212 17704 23252 17744
rect 23116 17620 23156 17660
rect 22924 17032 22964 17072
rect 23788 18460 23828 18500
rect 23980 18460 24020 18500
rect 23596 18040 23636 18080
rect 25228 18628 25268 18668
rect 26668 19132 26708 19172
rect 26572 18712 26612 18752
rect 24364 18376 24404 18416
rect 24172 18124 24212 18164
rect 25612 18544 25652 18584
rect 24556 18040 24596 18080
rect 25420 18040 25460 18080
rect 24172 17872 24212 17912
rect 26668 18544 26708 18584
rect 26956 20056 26996 20096
rect 27916 22072 27956 22112
rect 28204 22072 28244 22112
rect 27628 21736 27668 21776
rect 27628 20896 27668 20936
rect 27628 20224 27668 20264
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 28780 21904 28820 21944
rect 28012 21736 28052 21776
rect 28396 21652 28436 21692
rect 27820 21400 27860 21440
rect 28012 20812 28052 20852
rect 27916 20644 27956 20684
rect 26860 19888 26900 19928
rect 27340 19888 27380 19928
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 27724 20056 27764 20096
rect 27916 19468 27956 19508
rect 27628 19300 27668 19340
rect 27052 18712 27092 18752
rect 26956 18544 26996 18584
rect 26860 18376 26900 18416
rect 26476 18124 26516 18164
rect 26380 17788 26420 17828
rect 25516 17620 25556 17660
rect 25516 17368 25556 17408
rect 26764 17536 26804 17576
rect 24556 17032 24596 17072
rect 26476 17032 26516 17072
rect 27052 18376 27092 18416
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 27436 17956 27476 17996
rect 26860 17368 26900 17408
rect 26860 17032 26900 17072
rect 27052 17032 27092 17072
rect 27724 17704 27764 17744
rect 27436 16780 27476 16820
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 29068 21568 29108 21608
rect 28876 20980 28916 21020
rect 28684 20812 28724 20852
rect 28492 20728 28532 20768
rect 28876 20728 28916 20768
rect 29068 20980 29108 21020
rect 28396 20644 28436 20684
rect 28780 20644 28820 20684
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 28204 20140 28244 20180
rect 28300 20056 28340 20096
rect 29068 20140 29108 20180
rect 29068 19972 29108 20012
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 29452 21904 29492 21944
rect 29644 22240 29684 22280
rect 30316 22240 30356 22280
rect 29548 21568 29588 21608
rect 30412 22072 30452 22112
rect 30796 23164 30836 23204
rect 30796 22660 30836 22700
rect 30988 23248 31028 23288
rect 30988 22576 31028 22616
rect 30892 22408 30932 22448
rect 30508 21736 30548 21776
rect 30892 21652 30932 21692
rect 29356 21064 29396 21104
rect 29260 20896 29300 20936
rect 30508 20896 30548 20936
rect 29260 20644 29300 20684
rect 29164 19888 29204 19928
rect 32524 24676 32564 24716
rect 31756 24256 31796 24296
rect 31468 23836 31508 23876
rect 31468 23668 31508 23708
rect 31276 23248 31316 23288
rect 31372 23164 31412 23204
rect 31660 23164 31700 23204
rect 31276 22240 31316 22280
rect 31180 21820 31220 21860
rect 31468 22408 31508 22448
rect 31468 21568 31508 21608
rect 31852 23920 31892 23960
rect 31948 23248 31988 23288
rect 31852 22660 31892 22700
rect 32332 24256 32372 24296
rect 32716 24592 32756 24632
rect 32140 23668 32180 23708
rect 33196 25264 33236 25304
rect 33292 24592 33332 24632
rect 33580 25852 33620 25892
rect 34348 26104 34388 26144
rect 34732 26104 34772 26144
rect 34636 25936 34676 25976
rect 34636 25096 34676 25136
rect 33580 24508 33620 24548
rect 34348 24508 34388 24548
rect 33196 24340 33236 24380
rect 33388 24340 33428 24380
rect 32332 23752 32372 23792
rect 32428 23668 32468 23708
rect 32332 23332 32372 23372
rect 32044 22576 32084 22616
rect 32428 23080 32468 23120
rect 32812 23920 32852 23960
rect 32716 23248 32756 23288
rect 32620 23164 32660 23204
rect 32044 22240 32084 22280
rect 31756 22072 31796 22112
rect 31372 21232 31412 21272
rect 31180 20896 31220 20936
rect 31180 20728 31220 20768
rect 31660 20980 31700 21020
rect 32044 21988 32084 22028
rect 32044 21820 32084 21860
rect 32524 21988 32564 22028
rect 32332 21736 32372 21776
rect 34444 24256 34484 24296
rect 33388 23668 33428 23708
rect 33196 23164 33236 23204
rect 32812 23080 32852 23120
rect 33004 23080 33044 23120
rect 33292 23080 33332 23120
rect 34348 23752 34388 23792
rect 34540 23920 34580 23960
rect 34540 23500 34580 23540
rect 34444 23416 34484 23456
rect 32716 22660 32756 22700
rect 31852 20812 31892 20852
rect 31756 20140 31796 20180
rect 31468 19972 31508 20012
rect 31084 19216 31124 19256
rect 31660 19048 31700 19088
rect 29068 18628 29108 18668
rect 29932 18628 29972 18668
rect 30604 18628 30644 18668
rect 28684 18544 28724 18584
rect 28012 18208 28052 18248
rect 28972 18544 29012 18584
rect 29260 18292 29300 18332
rect 28780 18124 28820 18164
rect 27916 18040 27956 18080
rect 29836 18376 29876 18416
rect 30220 18376 30260 18416
rect 29740 17872 29780 17912
rect 27916 17704 27956 17744
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 27820 17032 27860 17072
rect 29164 17200 29204 17240
rect 27532 16192 27572 16232
rect 21964 16108 22004 16148
rect 27436 16108 27476 16148
rect 27820 16108 27860 16148
rect 21580 15940 21620 15980
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 9004 15352 9044 15392
rect 7468 15184 7508 15224
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 7468 14680 7508 14720
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 5932 12328 5972 12368
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 7468 12328 7508 12368
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 7468 11740 7508 11780
rect 7372 11572 7412 11612
rect 7180 9724 7220 9764
rect 7180 8632 7220 8672
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 29644 16780 29684 16820
rect 29644 16192 29684 16232
rect 29740 15772 29780 15812
rect 30124 18292 30164 18332
rect 30220 17956 30260 17996
rect 30028 17620 30068 17660
rect 29932 17536 29972 17576
rect 30412 17620 30452 17660
rect 31276 18460 31316 18500
rect 31180 18292 31220 18332
rect 31276 17788 31316 17828
rect 31852 19048 31892 19088
rect 31852 18628 31892 18668
rect 32140 20812 32180 20852
rect 32044 20224 32084 20264
rect 31756 18124 31796 18164
rect 31660 17704 31700 17744
rect 31564 17536 31604 17576
rect 30508 17200 30548 17240
rect 30700 17032 30740 17072
rect 30988 15688 31028 15728
rect 29836 15436 29876 15476
rect 29932 14596 29972 14636
rect 31180 14680 31220 14720
rect 31372 14596 31412 14636
rect 31948 17368 31988 17408
rect 31948 17032 31988 17072
rect 32908 22072 32948 22112
rect 32428 21232 32468 21272
rect 32428 20980 32468 21020
rect 32236 19972 32276 20012
rect 32236 19804 32276 19844
rect 32140 19552 32180 19592
rect 33004 21568 33044 21608
rect 33004 20896 33044 20936
rect 32908 20056 32948 20096
rect 32716 19804 32756 19844
rect 32140 18544 32180 18584
rect 32332 18544 32372 18584
rect 32140 18208 32180 18248
rect 32236 17704 32276 17744
rect 31756 15268 31796 15308
rect 31948 15520 31988 15560
rect 32044 15268 32084 15308
rect 32140 14512 32180 14552
rect 32524 18460 32564 18500
rect 32812 19720 32852 19760
rect 32908 19636 32948 19676
rect 34924 26356 34964 26396
rect 35020 26188 35060 26228
rect 35404 26356 35444 26396
rect 35212 25768 35252 25808
rect 35020 25516 35060 25556
rect 35788 25768 35828 25808
rect 35692 25516 35732 25556
rect 35500 25348 35540 25388
rect 35884 25348 35924 25388
rect 35692 25264 35732 25304
rect 35884 25096 35924 25136
rect 36364 25264 36404 25304
rect 35980 24760 36020 24800
rect 35212 24592 35252 24632
rect 35116 24004 35156 24044
rect 34828 23584 34868 23624
rect 35500 24088 35540 24128
rect 35500 23668 35540 23708
rect 35212 23248 35252 23288
rect 35884 24004 35924 24044
rect 35788 23500 35828 23540
rect 35884 23080 35924 23120
rect 36460 25096 36500 25136
rect 36076 23416 36116 23456
rect 36172 23332 36212 23372
rect 36364 23752 36404 23792
rect 36364 23164 36404 23204
rect 36076 23080 36116 23120
rect 36268 23080 36308 23120
rect 34924 22576 34964 22616
rect 35596 22408 35636 22448
rect 34924 21820 34964 21860
rect 35788 21736 35828 21776
rect 34636 21064 34676 21104
rect 33580 20728 33620 20768
rect 33196 19804 33236 19844
rect 33100 19720 33140 19760
rect 33196 19552 33236 19592
rect 32812 18544 32852 18584
rect 32524 17536 32564 17576
rect 33004 17368 33044 17408
rect 32812 17284 32852 17324
rect 32524 16192 32564 16232
rect 32332 15604 32372 15644
rect 32332 14512 32372 14552
rect 32236 14176 32276 14216
rect 32332 14092 32372 14132
rect 31852 14008 31892 14048
rect 31660 13420 31700 13460
rect 31852 13168 31892 13208
rect 32428 13420 32468 13460
rect 32908 15772 32948 15812
rect 32812 15604 32852 15644
rect 33292 18796 33332 18836
rect 33388 18712 33428 18752
rect 33292 18544 33332 18584
rect 36172 22408 36212 22448
rect 36268 21736 36308 21776
rect 36172 21568 36212 21608
rect 36748 25936 36788 25976
rect 36652 24760 36692 24800
rect 36556 23836 36596 23876
rect 38092 26356 38132 26396
rect 38092 26020 38132 26060
rect 37228 25852 37268 25892
rect 36940 25264 36980 25304
rect 38092 25600 38132 25640
rect 38476 25264 38516 25304
rect 36844 25096 36884 25136
rect 37516 24760 37556 24800
rect 37708 24676 37748 24716
rect 36748 24424 36788 24464
rect 36940 23248 36980 23288
rect 36460 22912 36500 22952
rect 36748 23080 36788 23120
rect 37324 23752 37364 23792
rect 37228 23584 37268 23624
rect 37132 23248 37172 23288
rect 37036 23080 37076 23120
rect 37228 23164 37268 23204
rect 36652 22408 36692 22448
rect 36844 22408 36884 22448
rect 34636 20392 34676 20432
rect 35212 20392 35252 20432
rect 34828 20140 34868 20180
rect 35020 20140 35060 20180
rect 34732 20056 34772 20096
rect 34924 20056 34964 20096
rect 34828 19972 34868 20012
rect 35020 19888 35060 19928
rect 37132 20896 37172 20936
rect 36652 20728 36692 20768
rect 36268 20056 36308 20096
rect 33484 18544 33524 18584
rect 33676 18544 33716 18584
rect 34828 18628 34868 18668
rect 35596 18628 35636 18668
rect 35788 18628 35828 18668
rect 34252 18544 34292 18584
rect 33484 18208 33524 18248
rect 33292 17704 33332 17744
rect 33580 18124 33620 18164
rect 34156 17704 34196 17744
rect 33292 17368 33332 17408
rect 33964 17032 34004 17072
rect 34540 17032 34580 17072
rect 34348 16864 34388 16904
rect 33484 16360 33524 16400
rect 33964 16696 34004 16736
rect 33676 16360 33716 16400
rect 33580 16276 33620 16316
rect 33004 15520 33044 15560
rect 35500 18544 35540 18584
rect 35404 18292 35444 18332
rect 36172 18628 36212 18668
rect 36460 18628 36500 18668
rect 36844 18628 36884 18668
rect 35692 18460 35732 18500
rect 36172 17200 36212 17240
rect 34732 16192 34772 16232
rect 34924 16108 34964 16148
rect 35980 16108 36020 16148
rect 33964 15856 34004 15896
rect 34636 15856 34676 15896
rect 33484 15772 33524 15812
rect 33868 15688 33908 15728
rect 34636 15604 34676 15644
rect 33388 15436 33428 15476
rect 34444 15520 34484 15560
rect 33004 15268 33044 15308
rect 33004 14764 33044 14804
rect 32716 14176 32756 14216
rect 32716 13504 32756 13544
rect 32812 13420 32852 13460
rect 33004 14176 33044 14216
rect 35116 15352 35156 15392
rect 34252 14680 34292 14720
rect 34828 14176 34868 14216
rect 35596 14848 35636 14888
rect 35500 14764 35540 14804
rect 35212 14680 35252 14720
rect 34924 12580 34964 12620
rect 33868 11908 33908 11948
rect 34828 11908 34868 11948
rect 34828 11656 34868 11696
rect 35116 13000 35156 13040
rect 35404 14176 35444 14216
rect 35404 13252 35444 13292
rect 35020 12160 35060 12200
rect 35308 11656 35348 11696
rect 34924 11572 34964 11612
rect 36556 17704 36596 17744
rect 36844 17704 36884 17744
rect 37036 19216 37076 19256
rect 36940 17200 36980 17240
rect 37228 19972 37268 20012
rect 37228 19048 37268 19088
rect 37132 17284 37172 17324
rect 37420 20728 37460 20768
rect 38092 23668 38132 23708
rect 37900 23332 37940 23372
rect 37804 23164 37844 23204
rect 38284 23164 38324 23204
rect 37996 22912 38036 22952
rect 38188 22408 38228 22448
rect 38476 22492 38516 22532
rect 55372 37360 55412 37400
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 49132 36016 49172 36056
rect 50476 36016 50516 36056
rect 43948 35932 43988 35972
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 49612 35596 49652 35636
rect 45964 34504 46004 34544
rect 46540 34504 46580 34544
rect 46828 34504 46868 34544
rect 49228 34504 49268 34544
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43180 33244 43220 33284
rect 43948 33244 43988 33284
rect 42124 33160 42164 33200
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 40972 31648 41012 31688
rect 41836 31648 41876 31688
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 40588 30556 40628 30596
rect 41164 30556 41204 30596
rect 40108 30388 40148 30428
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 40588 30136 40628 30176
rect 39532 30052 39572 30092
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 40012 29968 40052 30008
rect 40780 29968 40820 30008
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 41932 31144 41972 31184
rect 41836 30304 41876 30344
rect 40972 30220 41012 30260
rect 41356 30220 41396 30260
rect 41836 30136 41876 30176
rect 41644 30052 41684 30092
rect 40876 29128 40916 29168
rect 40204 28960 40244 29000
rect 40108 28708 40148 28748
rect 39724 28288 39764 28328
rect 38860 26020 38900 26060
rect 39724 27280 39764 27320
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 39148 27028 39188 27068
rect 39916 27028 39956 27068
rect 39340 26860 39380 26900
rect 39532 26860 39572 26900
rect 39052 26692 39092 26732
rect 40012 26776 40052 26816
rect 40492 28288 40532 28328
rect 41452 29800 41492 29840
rect 42028 30892 42068 30932
rect 41356 29716 41396 29756
rect 41356 29128 41396 29168
rect 41356 28876 41396 28916
rect 41260 28792 41300 28832
rect 41068 28540 41108 28580
rect 45868 33076 45908 33116
rect 42220 32908 42260 32948
rect 42796 32908 42836 32948
rect 42316 31564 42356 31604
rect 42220 30808 42260 30848
rect 42124 30556 42164 30596
rect 42508 31984 42548 32024
rect 42508 31648 42548 31688
rect 42508 31144 42548 31184
rect 42508 30808 42548 30848
rect 42412 30556 42452 30596
rect 42124 29716 42164 29756
rect 41644 29128 41684 29168
rect 41548 28876 41588 28916
rect 41452 28540 41492 28580
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 40492 27700 40532 27740
rect 40204 27532 40244 27572
rect 40204 27028 40244 27068
rect 39052 26272 39092 26312
rect 39436 26104 39476 26144
rect 39340 25936 39380 25976
rect 39244 25852 39284 25892
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 41356 28120 41396 28160
rect 41068 27532 41108 27572
rect 40588 27196 40628 27236
rect 41068 27196 41108 27236
rect 40876 27028 40916 27068
rect 40972 26860 41012 26900
rect 40492 26608 40532 26648
rect 40780 26608 40820 26648
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 40780 26440 40820 26480
rect 40588 26272 40628 26312
rect 40300 26104 40340 26144
rect 40204 25936 40244 25976
rect 38956 25264 38996 25304
rect 39916 25180 39956 25220
rect 40396 26020 40436 26060
rect 40876 26020 40916 26060
rect 41740 28960 41780 29000
rect 41740 28624 41780 28664
rect 42028 29128 42068 29168
rect 42124 29044 42164 29084
rect 41836 28540 41876 28580
rect 41932 28456 41972 28496
rect 41548 27784 41588 27824
rect 41644 27364 41684 27404
rect 42316 29800 42356 29840
rect 42316 29128 42356 29168
rect 43084 31564 43124 31604
rect 42988 31396 43028 31436
rect 42988 31144 43028 31184
rect 43372 30976 43412 31016
rect 43756 31312 43796 31352
rect 43276 30556 43316 30596
rect 43084 30472 43124 30512
rect 42796 30388 42836 30428
rect 42604 30304 42644 30344
rect 42412 28708 42452 28748
rect 42316 28456 42356 28496
rect 41452 26860 41492 26900
rect 41068 26104 41108 26144
rect 40108 25096 40148 25136
rect 39052 24508 39092 24548
rect 39532 24424 39572 24464
rect 39244 24340 39284 24380
rect 39820 24508 39860 24548
rect 39628 24256 39668 24296
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 38860 23668 38900 23708
rect 39052 23500 39092 23540
rect 38956 23416 38996 23456
rect 38860 23248 38900 23288
rect 40492 25516 40532 25556
rect 40780 25852 40820 25892
rect 41548 26608 41588 26648
rect 42028 26272 42068 26312
rect 41452 26104 41492 26144
rect 41644 26104 41684 26144
rect 40876 25516 40916 25556
rect 40684 25348 40724 25388
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 40492 24760 40532 24800
rect 40396 24592 40436 24632
rect 40108 24340 40148 24380
rect 39340 23164 39380 23204
rect 39724 23080 39764 23120
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 39052 22492 39092 22532
rect 39244 22240 39284 22280
rect 38572 21316 38612 21356
rect 38188 20392 38228 20432
rect 37804 20056 37844 20096
rect 37996 20056 38036 20096
rect 39244 21484 39284 21524
rect 39148 21400 39188 21440
rect 39052 21316 39092 21356
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 40012 23080 40052 23120
rect 39916 21400 39956 21440
rect 40684 24592 40724 24632
rect 40876 24760 40916 24800
rect 40972 24592 41012 24632
rect 41068 24508 41108 24548
rect 40876 24424 40916 24464
rect 41164 24256 41204 24296
rect 41164 23920 41204 23960
rect 40396 23668 40436 23708
rect 40876 23668 40916 23708
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 40204 22828 40244 22868
rect 40396 22324 40436 22364
rect 40588 22324 40628 22364
rect 41356 24424 41396 24464
rect 40876 23248 40916 23288
rect 41260 23332 41300 23372
rect 40780 22240 40820 22280
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 41068 21736 41108 21776
rect 41356 23248 41396 23288
rect 41452 22912 41492 22952
rect 41548 22660 41588 22700
rect 41260 21736 41300 21776
rect 41740 25852 41780 25892
rect 42796 29968 42836 30008
rect 42892 29128 42932 29168
rect 42796 27448 42836 27488
rect 43948 30976 43988 31016
rect 43948 30472 43988 30512
rect 44236 30640 44276 30680
rect 44140 30136 44180 30176
rect 44044 30052 44084 30092
rect 45964 32740 46004 32780
rect 46252 32320 46292 32360
rect 45676 32068 45716 32108
rect 45004 31648 45044 31688
rect 45100 30892 45140 30932
rect 45004 30724 45044 30764
rect 44908 30640 44948 30680
rect 44524 30220 44564 30260
rect 45100 30304 45140 30344
rect 44908 30052 44948 30092
rect 44524 29800 44564 29840
rect 44812 29800 44852 29840
rect 43852 29128 43892 29168
rect 46060 31564 46100 31604
rect 46156 31312 46196 31352
rect 45676 30556 45716 30596
rect 45292 30388 45332 30428
rect 45676 29548 45716 29588
rect 43564 28960 43604 29000
rect 43468 28792 43508 28832
rect 44620 28540 44660 28580
rect 43564 28288 43604 28328
rect 44332 27784 44372 27824
rect 43180 27616 43220 27656
rect 45100 28960 45140 29000
rect 46060 30640 46100 30680
rect 45964 30388 46004 30428
rect 46732 33160 46772 33200
rect 46348 30892 46388 30932
rect 46828 33076 46868 33116
rect 46924 32824 46964 32864
rect 46540 32404 46580 32444
rect 46636 32320 46676 32360
rect 47212 32740 47252 32780
rect 47308 32404 47348 32444
rect 46540 32068 46580 32108
rect 46444 30724 46484 30764
rect 46156 30136 46196 30176
rect 45964 30052 46004 30092
rect 46540 30556 46580 30596
rect 46348 30388 46388 30428
rect 46060 29380 46100 29420
rect 45388 28540 45428 28580
rect 46348 29380 46388 29420
rect 47116 32152 47156 32192
rect 48460 34336 48500 34376
rect 49228 34084 49268 34124
rect 48556 33160 48596 33200
rect 47596 33076 47636 33116
rect 48076 32992 48116 33032
rect 47404 32152 47444 32192
rect 47212 31312 47252 31352
rect 47692 32824 47732 32864
rect 48268 32824 48308 32864
rect 48268 32404 48308 32444
rect 48460 32152 48500 32192
rect 48076 31144 48116 31184
rect 47500 30640 47540 30680
rect 48652 32992 48692 33032
rect 49132 33664 49172 33704
rect 49036 33076 49076 33116
rect 48940 32992 48980 33032
rect 48844 32824 48884 32864
rect 48844 31732 48884 31772
rect 48652 31312 48692 31352
rect 48844 30976 48884 31016
rect 47116 30556 47156 30596
rect 45772 28372 45812 28412
rect 44908 28288 44948 28328
rect 45100 28288 45140 28328
rect 44812 28036 44852 28076
rect 44716 27952 44756 27992
rect 44620 27868 44660 27908
rect 44524 27280 44564 27320
rect 44716 27616 44756 27656
rect 45100 27616 45140 27656
rect 44620 27112 44660 27152
rect 43084 26776 43124 26816
rect 43564 26776 43604 26816
rect 41740 23416 41780 23456
rect 41836 23248 41876 23288
rect 42316 24592 42356 24632
rect 42124 23080 42164 23120
rect 41644 22324 41684 22364
rect 41548 21652 41588 21692
rect 40108 21484 40148 21524
rect 40972 20560 41012 20600
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 39628 20140 39668 20180
rect 40972 20140 41012 20180
rect 37612 19804 37652 19844
rect 38380 19804 38420 19844
rect 38668 19804 38708 19844
rect 37516 19468 37556 19508
rect 38188 19216 38228 19256
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 41260 21568 41300 21608
rect 41164 20560 41204 20600
rect 41164 20224 41204 20264
rect 42028 22912 42068 22952
rect 42412 22996 42452 23036
rect 42604 22828 42644 22868
rect 42124 22240 42164 22280
rect 42316 22240 42356 22280
rect 42316 21652 42356 21692
rect 42412 21484 42452 21524
rect 42316 21400 42356 21440
rect 41740 20728 41780 20768
rect 41644 20476 41684 20516
rect 41452 20140 41492 20180
rect 39052 19468 39092 19508
rect 41932 20224 41972 20264
rect 39148 19384 39188 19424
rect 38668 19048 38708 19088
rect 38380 18964 38420 19004
rect 37420 18544 37460 18584
rect 37420 17200 37460 17240
rect 36652 16864 36692 16904
rect 36268 16192 36308 16232
rect 36460 16192 36500 16232
rect 36172 16024 36212 16064
rect 36172 15772 36212 15812
rect 37132 16864 37172 16904
rect 37036 16780 37076 16820
rect 37036 16108 37076 16148
rect 36076 15520 36116 15560
rect 36076 14764 36116 14804
rect 36844 15520 36884 15560
rect 36268 15436 36308 15476
rect 36940 14848 36980 14888
rect 36844 14680 36884 14720
rect 36172 13840 36212 13880
rect 36076 13252 36116 13292
rect 36268 13420 36308 13460
rect 36268 13252 36308 13292
rect 37324 16444 37364 16484
rect 38572 17872 38612 17912
rect 38572 17032 38612 17072
rect 37708 16780 37748 16820
rect 37420 16360 37460 16400
rect 37996 16444 38036 16484
rect 37804 16192 37844 16232
rect 37996 16192 38036 16232
rect 37420 15856 37460 15896
rect 37516 15520 37556 15560
rect 37228 14008 37268 14048
rect 37804 14176 37844 14216
rect 37420 14092 37460 14132
rect 37804 14008 37844 14048
rect 37324 13840 37364 13880
rect 37132 13504 37172 13544
rect 36556 13168 36596 13208
rect 36076 12496 36116 12536
rect 35596 11656 35636 11696
rect 36076 11656 36116 11696
rect 36268 12496 36308 12536
rect 36364 12412 36404 12452
rect 37036 13168 37076 13208
rect 36844 13084 36884 13124
rect 36748 12496 36788 12536
rect 36652 12160 36692 12200
rect 37132 12664 37172 12704
rect 36844 11572 36884 11612
rect 35500 11404 35540 11444
rect 35404 10984 35444 11024
rect 36460 11488 36500 11528
rect 37036 11404 37076 11444
rect 36940 10984 36980 11024
rect 37132 10984 37172 11024
rect 36172 10816 36212 10856
rect 36748 10816 36788 10856
rect 38188 14932 38228 14972
rect 38092 14680 38132 14720
rect 38572 14680 38612 14720
rect 38380 14176 38420 14216
rect 38572 14092 38612 14132
rect 38092 13840 38132 13880
rect 38476 13924 38516 13964
rect 38284 13000 38324 13040
rect 38188 12496 38228 12536
rect 37996 11572 38036 11612
rect 38188 11488 38228 11528
rect 38956 19216 38996 19256
rect 38860 18628 38900 18668
rect 38860 13924 38900 13964
rect 38860 13168 38900 13208
rect 39724 19216 39764 19256
rect 39436 18964 39476 19004
rect 40684 19384 40724 19424
rect 40300 19300 40340 19340
rect 41260 19300 41300 19340
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 40972 18628 41012 18668
rect 39820 17704 39860 17744
rect 40204 18208 40244 18248
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 40012 17116 40052 17156
rect 39724 17032 39764 17072
rect 40876 16864 40916 16904
rect 39724 16780 39764 16820
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 39916 16612 39956 16652
rect 39628 16192 39668 16232
rect 39148 15520 39188 15560
rect 39244 15352 39284 15392
rect 39628 15604 39668 15644
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 39436 14932 39476 14972
rect 39628 14596 39668 14636
rect 40108 16192 40148 16232
rect 40012 15940 40052 15980
rect 40012 15772 40052 15812
rect 40780 15940 40820 15980
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 40204 15520 40244 15560
rect 40588 15520 40628 15560
rect 41164 18880 41204 18920
rect 41644 19048 41684 19088
rect 41452 18712 41492 18752
rect 41836 19300 41876 19340
rect 42124 20140 42164 20180
rect 41548 18040 41588 18080
rect 41068 17956 41108 17996
rect 41068 17452 41108 17492
rect 41068 17284 41108 17324
rect 41548 17452 41588 17492
rect 41356 16864 41396 16904
rect 41260 16780 41300 16820
rect 40012 14512 40052 14552
rect 39340 14260 39380 14300
rect 39148 14092 39188 14132
rect 39820 14176 39860 14216
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 41068 14344 41108 14384
rect 39244 13924 39284 13964
rect 40108 13840 40148 13880
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 40300 13420 40340 13460
rect 41164 14260 41204 14300
rect 44140 26608 44180 26648
rect 43852 25600 43892 25640
rect 44044 25600 44084 25640
rect 44908 27280 44948 27320
rect 44908 26020 44948 26060
rect 44332 25516 44372 25556
rect 44236 25432 44276 25472
rect 44620 25348 44660 25388
rect 44332 25264 44372 25304
rect 44428 24592 44468 24632
rect 44812 25852 44852 25892
rect 43276 24508 43316 24548
rect 43756 24424 43796 24464
rect 43276 23500 43316 23540
rect 44236 24340 44276 24380
rect 43852 24256 43892 24296
rect 43756 23248 43796 23288
rect 44044 24172 44084 24212
rect 43948 23752 43988 23792
rect 44140 23920 44180 23960
rect 44332 24172 44372 24212
rect 42988 22828 43028 22868
rect 43180 22744 43220 22784
rect 43468 22660 43508 22700
rect 43468 22492 43508 22532
rect 43084 22408 43124 22448
rect 42988 22324 43028 22364
rect 43564 22240 43604 22280
rect 42988 21820 43028 21860
rect 42412 20728 42452 20768
rect 42892 19972 42932 20012
rect 42508 19216 42548 19256
rect 42700 19216 42740 19256
rect 42124 18796 42164 18836
rect 42604 18628 42644 18668
rect 42028 18124 42068 18164
rect 42028 17956 42068 17996
rect 41932 17704 41972 17744
rect 41932 16948 41972 16988
rect 41836 16864 41876 16904
rect 42220 18376 42260 18416
rect 42892 19048 42932 19088
rect 42796 18712 42836 18752
rect 42412 18376 42452 18416
rect 42316 17956 42356 17996
rect 42124 17704 42164 17744
rect 42892 18208 42932 18248
rect 43660 20812 43700 20852
rect 44140 22912 44180 22952
rect 45868 28288 45908 28328
rect 45484 27952 45524 27992
rect 45676 27952 45716 27992
rect 45388 26104 45428 26144
rect 45292 25348 45332 25388
rect 45004 25264 45044 25304
rect 45292 25180 45332 25220
rect 44524 24172 44564 24212
rect 44908 24424 44948 24464
rect 44716 24340 44756 24380
rect 44620 23920 44660 23960
rect 44428 23752 44468 23792
rect 44620 23752 44660 23792
rect 44620 23248 44660 23288
rect 45100 24424 45140 24464
rect 45196 24340 45236 24380
rect 45100 23416 45140 23456
rect 44812 23332 44852 23372
rect 45004 23332 45044 23372
rect 44332 21400 44372 21440
rect 44620 20728 44660 20768
rect 45484 24340 45524 24380
rect 45388 24004 45428 24044
rect 45580 23080 45620 23120
rect 46060 28036 46100 28076
rect 46444 28288 46484 28328
rect 46636 28288 46676 28328
rect 46060 26356 46100 26396
rect 45964 26104 46004 26144
rect 46732 28204 46772 28244
rect 46636 28120 46676 28160
rect 46732 27952 46772 27992
rect 46540 27532 46580 27572
rect 48844 30472 48884 30512
rect 47788 30136 47828 30176
rect 49132 32068 49172 32108
rect 49036 31816 49076 31856
rect 48940 29884 48980 29924
rect 47788 29800 47828 29840
rect 48940 29380 48980 29420
rect 47308 28204 47348 28244
rect 46828 26776 46868 26816
rect 47404 27700 47444 27740
rect 47308 26776 47348 26816
rect 48844 28120 48884 28160
rect 47596 28036 47636 28076
rect 47692 27700 47732 27740
rect 47980 27616 48020 27656
rect 48652 27616 48692 27656
rect 47788 27532 47828 27572
rect 47020 26188 47060 26228
rect 46444 26020 46484 26060
rect 46348 25936 46388 25976
rect 46252 25852 46292 25892
rect 46540 25852 46580 25892
rect 46060 25768 46100 25808
rect 46348 25432 46388 25472
rect 46444 25264 46484 25304
rect 46732 25852 46772 25892
rect 46732 25096 46772 25136
rect 46828 25012 46868 25052
rect 47788 26104 47828 26144
rect 48844 26188 48884 26228
rect 49516 34336 49556 34376
rect 49228 31732 49268 31772
rect 50956 35932 50996 35972
rect 50476 35008 50516 35048
rect 50380 34672 50420 34712
rect 50092 34084 50132 34124
rect 49612 32152 49652 32192
rect 49420 32068 49460 32108
rect 49516 31480 49556 31520
rect 49324 31312 49364 31352
rect 49324 31144 49364 31184
rect 49420 30808 49460 30848
rect 49708 31480 49748 31520
rect 50092 32992 50132 33032
rect 49996 31732 50036 31772
rect 49420 30472 49460 30512
rect 49324 30220 49364 30260
rect 49228 29800 49268 29840
rect 49900 30724 49940 30764
rect 50476 34336 50516 34376
rect 51436 35848 51476 35888
rect 51436 35176 51476 35216
rect 51628 35260 51668 35300
rect 52780 35848 52820 35888
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 51532 35092 51572 35132
rect 51340 35008 51380 35048
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 51148 34588 51188 34628
rect 51532 34588 51572 34628
rect 50572 33076 50612 33116
rect 51244 34504 51284 34544
rect 51724 34672 51764 34712
rect 52108 35092 52148 35132
rect 52300 35176 52340 35216
rect 53260 35596 53300 35636
rect 54412 35596 54452 35636
rect 55660 37360 55700 37400
rect 55660 37192 55700 37232
rect 55564 36772 55604 36812
rect 57292 38032 57332 38072
rect 57196 37360 57236 37400
rect 57484 37276 57524 37316
rect 56716 37192 56756 37232
rect 55756 36856 55796 36896
rect 56236 36604 56276 36644
rect 55468 35764 55508 35804
rect 55180 35344 55220 35384
rect 54412 35260 54452 35300
rect 54796 35260 54836 35300
rect 55276 35260 55316 35300
rect 52780 34672 52820 34712
rect 52204 34504 52244 34544
rect 51820 34336 51860 34376
rect 50956 33664 50996 33704
rect 50668 32992 50708 33032
rect 50860 32824 50900 32864
rect 52396 34336 52436 34376
rect 52492 34168 52532 34208
rect 52204 34084 52244 34124
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 52204 33748 52244 33788
rect 53644 34168 53684 34208
rect 51532 33412 51572 33452
rect 51820 33412 51860 33452
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 51148 32992 51188 33032
rect 50572 32656 50612 32696
rect 50572 31984 50612 32024
rect 50668 31732 50708 31772
rect 51148 32824 51188 32864
rect 51244 32656 51284 32696
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 51148 31312 51188 31352
rect 51628 31396 51668 31436
rect 50860 30808 50900 30848
rect 50380 30724 50420 30764
rect 51820 32740 51860 32780
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 53644 33580 53684 33620
rect 53740 33076 53780 33116
rect 53836 32824 53876 32864
rect 54124 34336 54164 34376
rect 54124 34084 54164 34124
rect 54028 33748 54068 33788
rect 52396 32152 52436 32192
rect 53452 32152 53492 32192
rect 54604 33916 54644 33956
rect 54604 33580 54644 33620
rect 54316 33244 54356 33284
rect 54604 33076 54644 33116
rect 55852 35680 55892 35720
rect 55564 35260 55604 35300
rect 55084 35176 55124 35216
rect 54988 34672 55028 34712
rect 55180 34756 55220 34796
rect 55084 34336 55124 34376
rect 55276 33916 55316 33956
rect 55084 33832 55124 33872
rect 54796 33412 54836 33452
rect 54892 33328 54932 33368
rect 54700 32488 54740 32528
rect 54892 32824 54932 32864
rect 55276 33496 55316 33536
rect 55180 32824 55220 32864
rect 55372 33328 55412 33368
rect 54988 32572 55028 32612
rect 51916 31396 51956 31436
rect 50284 30304 50324 30344
rect 49516 29884 49556 29924
rect 49708 29800 49748 29840
rect 49996 29800 50036 29840
rect 49900 29716 49940 29756
rect 50764 30640 50804 30680
rect 50764 30388 50804 30428
rect 50476 29800 50516 29840
rect 48940 26104 48980 26144
rect 49132 26104 49172 26144
rect 47404 25936 47444 25976
rect 47116 24844 47156 24884
rect 47500 25012 47540 25052
rect 47308 24760 47348 24800
rect 46828 24592 46868 24632
rect 46348 24508 46388 24548
rect 47212 24592 47252 24632
rect 47308 24508 47348 24548
rect 47116 24256 47156 24296
rect 46252 24172 46292 24212
rect 46924 24172 46964 24212
rect 46060 23752 46100 23792
rect 45868 23080 45908 23120
rect 46156 23584 46196 23624
rect 46540 23332 46580 23372
rect 46156 23109 46196 23120
rect 46156 23080 46196 23109
rect 44908 21568 44948 21608
rect 45292 22996 45332 23036
rect 45004 21400 45044 21440
rect 44908 20728 44948 20768
rect 45388 22240 45428 22280
rect 45292 21988 45332 22028
rect 46156 22660 46196 22700
rect 45580 21904 45620 21944
rect 45196 21652 45236 21692
rect 45388 21568 45428 21608
rect 45292 21484 45332 21524
rect 46060 21988 46100 22028
rect 45676 21316 45716 21356
rect 45484 20812 45524 20852
rect 43276 19972 43316 20012
rect 43276 19804 43316 19844
rect 43276 19300 43316 19340
rect 43180 18880 43220 18920
rect 43468 18712 43508 18752
rect 43084 18460 43124 18500
rect 43276 18376 43316 18416
rect 42700 17788 42740 17828
rect 42124 16948 42164 16988
rect 41740 16780 41780 16820
rect 41644 16024 41684 16064
rect 41452 14680 41492 14720
rect 41356 14428 41396 14468
rect 41356 14260 41396 14300
rect 41260 14176 41300 14216
rect 41068 13924 41108 13964
rect 39340 13084 39380 13124
rect 38956 12664 38996 12704
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 39532 12664 39572 12704
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 38860 11656 38900 11696
rect 38764 10984 38804 11024
rect 38860 10564 38900 10604
rect 38668 10060 38708 10100
rect 29164 9472 29204 9512
rect 40300 12496 40340 12536
rect 39148 11656 39188 11696
rect 39532 11656 39572 11696
rect 39340 11572 39380 11612
rect 39628 11488 39668 11528
rect 39436 10984 39476 11024
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 39148 10228 39188 10268
rect 40012 10732 40052 10772
rect 39244 10060 39284 10100
rect 39340 9640 39380 9680
rect 39436 9472 39476 9512
rect 40588 9976 40628 10016
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 40876 10060 40916 10100
rect 40108 9640 40148 9680
rect 40780 9640 40820 9680
rect 40684 9556 40724 9596
rect 40204 9472 40244 9512
rect 40588 9472 40628 9512
rect 42028 15604 42068 15644
rect 41548 13420 41588 13460
rect 41740 13168 41780 13208
rect 42220 15604 42260 15644
rect 42028 14680 42068 14720
rect 41932 13840 41972 13880
rect 41452 12580 41492 12620
rect 41740 12496 41780 12536
rect 41452 11740 41492 11780
rect 41836 12244 41876 12284
rect 42316 13840 42356 13880
rect 42604 16948 42644 16988
rect 42892 17704 42932 17744
rect 42796 17620 42836 17660
rect 42892 16864 42932 16904
rect 42508 16192 42548 16232
rect 42700 16612 42740 16652
rect 43180 17620 43220 17660
rect 43372 17284 43412 17324
rect 42892 16192 42932 16232
rect 43276 15856 43316 15896
rect 43084 15604 43124 15644
rect 45676 20728 45716 20768
rect 45964 21316 46004 21356
rect 46060 20728 46100 20768
rect 46252 22240 46292 22280
rect 46348 20728 46388 20768
rect 46732 23164 46772 23204
rect 46636 22240 46676 22280
rect 47692 23920 47732 23960
rect 48364 23920 48404 23960
rect 48556 24256 48596 24296
rect 47980 23584 48020 23624
rect 48844 24004 48884 24044
rect 48652 23248 48692 23288
rect 46732 20728 46772 20768
rect 44524 19972 44564 20012
rect 44140 19888 44180 19928
rect 43852 19804 43892 19844
rect 44812 20224 44852 20264
rect 44716 19888 44756 19928
rect 44332 19216 44372 19256
rect 43660 18544 43700 18584
rect 43756 18460 43796 18500
rect 43948 18628 43988 18668
rect 44044 18544 44084 18584
rect 44236 18544 44276 18584
rect 44236 18292 44276 18332
rect 43948 17788 43988 17828
rect 44140 17704 44180 17744
rect 44620 18880 44660 18920
rect 44524 18544 44564 18584
rect 44428 18376 44468 18416
rect 44620 18376 44660 18416
rect 44716 18040 44756 18080
rect 44044 16864 44084 16904
rect 43852 16696 43892 16736
rect 43660 15352 43700 15392
rect 44716 16864 44756 16904
rect 44524 16696 44564 16736
rect 44332 16024 44372 16064
rect 44524 16024 44564 16064
rect 44236 15352 44276 15392
rect 42604 14680 42644 14720
rect 42604 14176 42644 14216
rect 42796 14680 42836 14720
rect 43084 14680 43124 14720
rect 43372 14680 43412 14720
rect 42604 13336 42644 13376
rect 42316 12832 42356 12872
rect 42412 12496 42452 12536
rect 42316 12244 42356 12284
rect 42412 11992 42452 12032
rect 42124 11320 42164 11360
rect 41548 10816 41588 10856
rect 42124 11152 42164 11192
rect 42508 11152 42548 11192
rect 42028 10732 42068 10772
rect 42796 13168 42836 13208
rect 43180 14092 43220 14132
rect 43372 14092 43412 14132
rect 43564 14092 43604 14132
rect 43276 13420 43316 13460
rect 42700 13000 42740 13040
rect 43468 13672 43508 13712
rect 44332 14092 44372 14132
rect 43852 13672 43892 13712
rect 43660 13000 43700 13040
rect 42988 12832 43028 12872
rect 42508 10732 42548 10772
rect 42124 10396 42164 10436
rect 41740 10060 41780 10100
rect 42220 10060 42260 10100
rect 41836 9976 41876 10016
rect 41356 9556 41396 9596
rect 41740 9808 41780 9848
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 41548 9220 41588 9260
rect 41452 8632 41492 8672
rect 41932 9556 41972 9596
rect 42316 9892 42356 9932
rect 42796 9640 42836 9680
rect 42700 9472 42740 9512
rect 44428 13000 44468 13040
rect 43564 11656 43604 11696
rect 44332 11656 44372 11696
rect 43948 11236 43988 11276
rect 43468 11152 43508 11192
rect 43852 11152 43892 11192
rect 43084 10816 43124 10856
rect 43084 10144 43124 10184
rect 43468 10144 43508 10184
rect 45004 20140 45044 20180
rect 45196 20056 45236 20096
rect 45004 19216 45044 19256
rect 45100 18460 45140 18500
rect 44908 18040 44948 18080
rect 45100 16780 45140 16820
rect 45292 19972 45332 20012
rect 45580 18712 45620 18752
rect 45484 18628 45524 18668
rect 45484 18376 45524 18416
rect 45292 18124 45332 18164
rect 45196 15184 45236 15224
rect 45388 16864 45428 16904
rect 46636 19972 46676 20012
rect 46156 18712 46196 18752
rect 46156 18544 46196 18584
rect 46252 18376 46292 18416
rect 45868 18292 45908 18332
rect 45676 18040 45716 18080
rect 46444 18460 46484 18500
rect 45964 18124 46004 18164
rect 45868 17956 45908 17996
rect 46348 17956 46388 17996
rect 45964 17620 46004 17660
rect 46348 17620 46388 17660
rect 46540 18208 46580 18248
rect 46156 17536 46196 17576
rect 46444 17536 46484 17576
rect 47692 21316 47732 21356
rect 47212 20728 47252 20768
rect 47596 20728 47636 20768
rect 48556 22240 48596 22280
rect 48748 23164 48788 23204
rect 49228 25936 49268 25976
rect 49516 27532 49556 27572
rect 49516 26356 49556 26396
rect 49420 25684 49460 25724
rect 49804 28960 49844 29000
rect 50668 29800 50708 29840
rect 50572 29632 50612 29672
rect 51148 30724 51188 30764
rect 51724 30724 51764 30764
rect 51244 30388 51284 30428
rect 51820 30640 51860 30680
rect 51532 30556 51572 30596
rect 54412 32068 54452 32108
rect 53548 31984 53588 32024
rect 52108 31312 52148 31352
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 52108 30808 52148 30848
rect 51628 30472 51668 30512
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 51724 30388 51764 30428
rect 51724 30220 51764 30260
rect 51532 29632 51572 29672
rect 50380 28960 50420 29000
rect 49996 28708 50036 28748
rect 50188 28456 50228 28496
rect 49996 28288 50036 28328
rect 50956 28792 50996 28832
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 51340 28540 51380 28580
rect 51724 28456 51764 28496
rect 50476 28288 50516 28328
rect 50572 28204 50612 28244
rect 50764 28288 50804 28328
rect 50092 28120 50132 28160
rect 50668 28120 50708 28160
rect 50092 27616 50132 27656
rect 50572 27532 50612 27572
rect 50398 26944 50438 26984
rect 50284 26608 50324 26648
rect 49996 25684 50036 25724
rect 49228 23920 49268 23960
rect 49516 25012 49556 25052
rect 49516 24676 49556 24716
rect 50188 25264 50228 25304
rect 51244 28288 51284 28328
rect 50956 28204 50996 28244
rect 50764 26608 50804 26648
rect 51532 27952 51572 27992
rect 51628 27700 51668 27740
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 51436 26608 51476 26648
rect 51148 26272 51188 26312
rect 51820 27196 51860 27236
rect 52204 30556 52244 30596
rect 52108 30220 52148 30260
rect 53452 31312 53492 31352
rect 54028 31312 54068 31352
rect 54892 32068 54932 32108
rect 54796 31900 54836 31940
rect 54700 30640 54740 30680
rect 52300 30472 52340 30512
rect 52780 30472 52820 30512
rect 54508 30472 54548 30512
rect 52492 30136 52532 30176
rect 52012 28120 52052 28160
rect 52012 27952 52052 27992
rect 52012 27700 52052 27740
rect 54796 29884 54836 29924
rect 52492 29800 52532 29840
rect 54124 29800 54164 29840
rect 53644 29632 53684 29672
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 52300 29044 52340 29084
rect 54316 29632 54356 29672
rect 54124 29128 54164 29168
rect 53260 29044 53300 29084
rect 52876 28456 52916 28496
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 52108 27196 52148 27236
rect 51532 26188 51572 26228
rect 50668 26104 50708 26144
rect 50572 25432 50612 25472
rect 50668 25264 50708 25304
rect 50476 24676 50516 24716
rect 49804 24340 49844 24380
rect 50188 24340 50228 24380
rect 50380 24340 50420 24380
rect 49900 23920 49940 23960
rect 49804 23248 49844 23288
rect 49708 23080 49748 23120
rect 49996 23752 50036 23792
rect 49900 23164 49940 23204
rect 49036 22324 49076 22364
rect 48940 22240 48980 22280
rect 48364 21484 48404 21524
rect 49228 22072 49268 22112
rect 50956 25936 50996 25976
rect 51244 25852 51284 25892
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 50956 24844 50996 24884
rect 50860 24340 50900 24380
rect 50764 23920 50804 23960
rect 50572 23752 50612 23792
rect 50380 23332 50420 23372
rect 50668 23584 50708 23624
rect 51340 25096 51380 25136
rect 51148 24592 51188 24632
rect 51724 26104 51764 26144
rect 53164 28120 53204 28160
rect 52972 26776 53012 26816
rect 52204 26608 52244 26648
rect 52012 26524 52052 26564
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 52108 26272 52148 26312
rect 52012 26188 52052 26228
rect 52492 26188 52532 26228
rect 51820 25936 51860 25976
rect 51724 25852 51764 25892
rect 51724 25432 51764 25472
rect 51820 25264 51860 25304
rect 52012 25180 52052 25220
rect 51916 25096 51956 25136
rect 51820 24928 51860 24968
rect 51628 24592 51668 24632
rect 51052 23920 51092 23960
rect 51052 23752 51092 23792
rect 50769 23584 50809 23624
rect 50572 23416 50612 23456
rect 50476 23164 50516 23204
rect 50188 22996 50228 23036
rect 50764 23248 50804 23288
rect 50668 23164 50708 23204
rect 50284 22156 50324 22196
rect 49036 21568 49076 21608
rect 50380 21988 50420 22028
rect 49516 21904 49556 21944
rect 49612 21568 49652 21608
rect 48844 21316 48884 21356
rect 48556 20980 48596 21020
rect 50380 21652 50420 21692
rect 50092 20980 50132 21020
rect 48940 20728 48980 20768
rect 51244 23584 51284 23624
rect 51052 23248 51092 23288
rect 51436 23248 51476 23288
rect 51340 23080 51380 23120
rect 50860 22492 50900 22532
rect 50860 22156 50900 22196
rect 50764 22072 50804 22112
rect 50764 21736 50804 21776
rect 51724 23584 51764 23624
rect 51724 23416 51764 23456
rect 51820 23332 51860 23372
rect 51820 23164 51860 23204
rect 51532 22996 51572 23036
rect 51820 22744 51860 22784
rect 51436 22240 51476 22280
rect 51148 21904 51188 21944
rect 51148 21736 51188 21776
rect 51052 21652 51092 21692
rect 50956 21568 50996 21608
rect 50860 20728 50900 20768
rect 51532 20728 51572 20768
rect 47596 20140 47636 20180
rect 47308 19804 47348 19844
rect 47020 19468 47060 19508
rect 47500 19804 47540 19844
rect 47404 18880 47444 18920
rect 47692 19804 47732 19844
rect 49324 19972 49364 20012
rect 46828 18628 46868 18668
rect 47020 18544 47060 18584
rect 47404 18544 47444 18584
rect 46924 18460 46964 18500
rect 46828 18376 46868 18416
rect 46732 17956 46772 17996
rect 46732 17536 46772 17576
rect 47500 18376 47540 18416
rect 46828 17284 46868 17324
rect 47692 18544 47732 18584
rect 45676 16948 45716 16988
rect 45868 16780 45908 16820
rect 45964 16528 46004 16568
rect 46252 16528 46292 16568
rect 45580 16108 45620 16148
rect 45484 16024 45524 16064
rect 45484 15688 45524 15728
rect 45580 15604 45620 15644
rect 45964 15856 46004 15896
rect 46252 16192 46292 16232
rect 46252 15604 46292 15644
rect 46060 15520 46100 15560
rect 47212 16864 47252 16904
rect 46444 15520 46484 15560
rect 48076 18628 48116 18668
rect 47980 18460 48020 18500
rect 48652 18544 48692 18584
rect 48460 18292 48500 18332
rect 48268 18124 48308 18164
rect 48460 17872 48500 17912
rect 48940 18880 48980 18920
rect 49132 19132 49172 19172
rect 49036 18712 49076 18752
rect 49228 18712 49268 18752
rect 51628 19972 51668 20012
rect 49612 19132 49652 19172
rect 50860 18796 50900 18836
rect 48940 18544 48980 18584
rect 48844 18460 48884 18500
rect 48748 18376 48788 18416
rect 48940 17872 48980 17912
rect 48748 17536 48788 17576
rect 47980 17368 48020 17408
rect 48940 17368 48980 17408
rect 48844 17284 48884 17324
rect 48268 17200 48308 17240
rect 48652 16948 48692 16988
rect 48268 16864 48308 16904
rect 48652 16192 48692 16232
rect 47404 15604 47444 15644
rect 45580 14932 45620 14972
rect 46156 14932 46196 14972
rect 45772 14764 45812 14804
rect 45484 13420 45524 13460
rect 44812 12664 44852 12704
rect 44716 12160 44756 12200
rect 44620 11992 44660 12032
rect 45868 14680 45908 14720
rect 46348 14680 46388 14720
rect 46252 14596 46292 14636
rect 46060 14344 46100 14384
rect 45868 14092 45908 14132
rect 46252 14092 46292 14132
rect 46156 14008 46196 14048
rect 46060 13336 46100 13376
rect 46252 13000 46292 13040
rect 45580 12244 45620 12284
rect 45484 11908 45524 11948
rect 44524 11824 44564 11864
rect 44908 11824 44948 11864
rect 45388 11656 45428 11696
rect 48076 15604 48116 15644
rect 47212 15352 47252 15392
rect 47980 15520 48020 15560
rect 47788 15352 47828 15392
rect 47308 14680 47348 14720
rect 46924 14512 46964 14552
rect 46540 14344 46580 14384
rect 47404 14344 47444 14384
rect 47596 14092 47636 14132
rect 46540 14008 46580 14048
rect 47500 14008 47540 14048
rect 47788 14008 47828 14048
rect 49132 17284 49172 17324
rect 49900 18544 49940 18584
rect 49516 18460 49556 18500
rect 49420 18292 49460 18332
rect 49900 18292 49940 18332
rect 49324 18208 49364 18248
rect 49420 17872 49460 17912
rect 49228 17200 49268 17240
rect 49228 16864 49268 16904
rect 49324 16780 49364 16820
rect 49132 15604 49172 15644
rect 48940 15268 48980 15308
rect 49228 14596 49268 14636
rect 48364 14512 48404 14552
rect 46636 13000 46676 13040
rect 47500 13252 47540 13292
rect 46828 12412 46868 12452
rect 46828 11992 46868 12032
rect 46540 11740 46580 11780
rect 47500 12832 47540 12872
rect 48076 13420 48116 13460
rect 47884 12664 47924 12704
rect 47020 12412 47060 12452
rect 46924 11656 46964 11696
rect 47116 11656 47156 11696
rect 48652 14344 48692 14384
rect 48460 13336 48500 13376
rect 49420 16192 49460 16232
rect 49900 17116 49940 17156
rect 49900 16780 49940 16820
rect 49900 15856 49940 15896
rect 50092 17704 50132 17744
rect 50572 18124 50612 18164
rect 50572 17872 50612 17912
rect 50476 17788 50516 17828
rect 50380 17704 50420 17744
rect 49036 14092 49076 14132
rect 49324 14092 49364 14132
rect 48460 13000 48500 13040
rect 48460 12748 48500 12788
rect 48556 12664 48596 12704
rect 48748 12664 48788 12704
rect 49516 13252 49556 13292
rect 49132 13084 49172 13124
rect 49420 13084 49460 13124
rect 49228 12664 49268 12704
rect 48268 11908 48308 11948
rect 48556 11824 48596 11864
rect 49132 11824 49172 11864
rect 48460 11656 48500 11696
rect 49324 12496 49364 12536
rect 49996 15520 50036 15560
rect 49996 15268 50036 15308
rect 49708 12832 49748 12872
rect 49708 12664 49748 12704
rect 49612 12496 49652 12536
rect 49612 12244 49652 12284
rect 49228 11656 49268 11696
rect 49420 11656 49460 11696
rect 49132 11488 49172 11528
rect 49804 11488 49844 11528
rect 46252 11236 46292 11276
rect 46540 11152 46580 11192
rect 46540 10816 46580 10856
rect 48076 11068 48116 11108
rect 46828 10396 46868 10436
rect 46252 10228 46292 10268
rect 43660 10060 43700 10100
rect 43276 9892 43316 9932
rect 43084 9640 43124 9680
rect 42988 9556 43028 9596
rect 42892 9472 42932 9512
rect 42412 9220 42452 9260
rect 41836 8716 41876 8756
rect 42796 8716 42836 8756
rect 41932 8632 41972 8672
rect 7660 8464 7700 8504
rect 6412 7960 6452 8000
rect 6316 5860 6356 5900
rect 6220 5608 6260 5648
rect 7468 7708 7508 7748
rect 7468 6532 7508 6572
rect 7468 6196 7508 6236
rect 6124 5188 6164 5228
rect 5932 5104 5972 5144
rect 4780 4180 4820 4220
rect 4876 4096 4916 4136
rect 5068 4096 5108 4136
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 4396 3508 4436 3548
rect 4876 3508 4916 3548
rect 3052 2584 3092 2624
rect 6508 5020 6548 5060
rect 6316 4096 6356 4136
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 43084 9304 43124 9344
rect 42988 8044 43028 8084
rect 44428 10060 44468 10100
rect 46348 10060 46388 10100
rect 43852 9472 43892 9512
rect 44524 9472 44564 9512
rect 45868 9472 45908 9512
rect 45388 9388 45428 9428
rect 44908 9220 44948 9260
rect 44236 8128 44276 8168
rect 44428 7960 44468 8000
rect 45004 8128 45044 8168
rect 45580 9304 45620 9344
rect 45484 8716 45524 8756
rect 44428 7792 44468 7832
rect 44812 7792 44852 7832
rect 43276 7708 43316 7748
rect 44236 7708 44276 7748
rect 45388 7708 45428 7748
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 46732 10060 46772 10100
rect 45964 9220 46004 9260
rect 46444 9220 46484 9260
rect 49324 10984 49364 11024
rect 47116 10396 47156 10436
rect 49132 10396 49172 10436
rect 48364 10312 48404 10352
rect 46924 9892 46964 9932
rect 46540 8716 46580 8756
rect 45484 6364 45524 6404
rect 45676 7960 45716 8000
rect 46924 8548 46964 8588
rect 47980 8716 48020 8756
rect 48172 8716 48212 8756
rect 47980 8548 48020 8588
rect 46732 7960 46772 8000
rect 47020 7960 47060 8000
rect 46828 7792 46868 7832
rect 47308 7960 47348 8000
rect 45580 6280 45620 6320
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 45676 5020 45716 5060
rect 47692 7876 47732 7916
rect 47500 7708 47540 7748
rect 47500 7372 47540 7412
rect 47116 6364 47156 6404
rect 47308 6364 47348 6404
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 7660 4264 7700 4304
rect 47884 7792 47924 7832
rect 47788 7372 47828 7412
rect 47980 7372 48020 7412
rect 47404 6280 47444 6320
rect 47404 5776 47444 5816
rect 47404 5608 47444 5648
rect 47596 5776 47636 5816
rect 47308 5020 47348 5060
rect 48844 10228 48884 10268
rect 48460 9472 48500 9512
rect 48460 8716 48500 8756
rect 48556 8548 48596 8588
rect 48268 8212 48308 8252
rect 48556 7960 48596 8000
rect 50476 16696 50516 16736
rect 50380 15352 50420 15392
rect 50668 17200 50708 17240
rect 51340 18376 51380 18416
rect 51340 17284 51380 17324
rect 51436 17200 51476 17240
rect 51340 17116 51380 17156
rect 50860 16612 50900 16652
rect 50764 15520 50804 15560
rect 51340 16864 51380 16904
rect 51724 18292 51764 18332
rect 52108 24928 52148 24968
rect 52684 25852 52724 25892
rect 52684 25264 52724 25304
rect 52876 25600 52916 25640
rect 52396 25180 52436 25220
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 52300 24592 52340 24632
rect 52204 24424 52244 24464
rect 52204 23920 52244 23960
rect 53293 27616 53333 27656
rect 53293 27448 53333 27488
rect 54220 27028 54260 27068
rect 53644 24592 53684 24632
rect 53164 24424 53204 24464
rect 54700 28792 54740 28832
rect 54604 28540 54644 28580
rect 54508 28456 54548 28496
rect 55180 32068 55220 32108
rect 56044 35848 56084 35888
rect 55660 33160 55700 33200
rect 55564 32488 55604 32528
rect 55468 31396 55508 31436
rect 55852 35092 55892 35132
rect 56044 35092 56084 35132
rect 56332 35764 56372 35804
rect 56620 35680 56660 35720
rect 57100 36856 57140 36896
rect 56812 35932 56852 35972
rect 56908 35848 56948 35888
rect 57292 36688 57332 36728
rect 57196 36604 57236 36644
rect 56428 34840 56468 34880
rect 55948 34504 55988 34544
rect 55948 34336 55988 34376
rect 56236 34336 56276 34376
rect 56524 34504 56564 34544
rect 56428 34420 56468 34460
rect 56332 34252 56372 34292
rect 55852 34000 55892 34040
rect 56236 34000 56276 34040
rect 56332 33244 56372 33284
rect 55756 31900 55796 31940
rect 55276 30976 55316 31016
rect 55084 30388 55124 30428
rect 54988 30220 55028 30260
rect 55180 29884 55220 29924
rect 54988 29800 55028 29840
rect 54988 29548 55028 29588
rect 54892 28708 54932 28748
rect 54892 28204 54932 28244
rect 54796 27616 54836 27656
rect 54892 27280 54932 27320
rect 54412 26692 54452 26732
rect 54700 26692 54740 26732
rect 54700 26272 54740 26312
rect 55084 29296 55124 29336
rect 55372 30724 55412 30764
rect 55660 30640 55700 30680
rect 57004 35176 57044 35216
rect 55948 30976 55988 31016
rect 55948 30808 55988 30848
rect 56140 30640 56180 30680
rect 56908 31312 56948 31352
rect 56620 31060 56660 31100
rect 56620 30724 56660 30764
rect 56236 30556 56276 30596
rect 55948 30304 55988 30344
rect 56332 30304 56372 30344
rect 56236 30220 56276 30260
rect 55468 29548 55508 29588
rect 55276 29296 55316 29336
rect 55276 28624 55316 28664
rect 55660 29548 55700 29588
rect 55468 28792 55508 28832
rect 55756 29296 55796 29336
rect 55564 28708 55604 28748
rect 55372 28120 55412 28160
rect 55468 27868 55508 27908
rect 55660 28288 55700 28328
rect 55948 28708 55988 28748
rect 56524 30556 56564 30596
rect 56428 29800 56468 29840
rect 57484 34924 57524 34964
rect 57580 33748 57620 33788
rect 57868 38116 57908 38156
rect 58060 37948 58100 37988
rect 58060 37276 58100 37316
rect 57964 34840 58004 34880
rect 58156 37192 58196 37232
rect 59404 38200 59444 38240
rect 59980 38032 60020 38072
rect 58348 37444 58388 37484
rect 58252 36856 58292 36896
rect 58540 36940 58580 36980
rect 58156 35176 58196 35216
rect 58156 34924 58196 34964
rect 58156 34588 58196 34628
rect 58060 34168 58100 34208
rect 57772 33916 57812 33956
rect 57772 33748 57812 33788
rect 57676 32992 57716 33032
rect 57772 32824 57812 32864
rect 58348 36688 58388 36728
rect 59788 37948 59828 37988
rect 58828 37360 58868 37400
rect 60460 38032 60500 38072
rect 60268 37444 60308 37484
rect 58732 37276 58772 37316
rect 58828 37192 58868 37232
rect 58636 36688 58676 36728
rect 59020 36856 59060 36896
rect 59788 36940 59828 36980
rect 59308 36856 59348 36896
rect 58444 35848 58484 35888
rect 58732 35848 58772 35888
rect 58348 34504 58388 34544
rect 58252 34336 58292 34376
rect 58828 34252 58868 34292
rect 58444 34168 58484 34208
rect 58348 33916 58388 33956
rect 59116 34588 59156 34628
rect 60364 37360 60404 37400
rect 61132 37948 61172 37988
rect 59788 34504 59828 34544
rect 59596 34420 59636 34460
rect 59212 34336 59252 34376
rect 58540 33412 58580 33452
rect 58060 32572 58100 32612
rect 57388 31312 57428 31352
rect 58444 32824 58484 32864
rect 58924 33412 58964 33452
rect 58732 33244 58772 33284
rect 58348 32740 58388 32780
rect 58348 32236 58388 32276
rect 58156 30808 58196 30848
rect 57772 30724 57812 30764
rect 58732 32740 58772 32780
rect 59692 33664 59732 33704
rect 59116 33076 59156 33116
rect 59404 33076 59444 33116
rect 58636 32488 58676 32528
rect 59020 32488 59060 32528
rect 58828 32320 58868 32360
rect 58444 32068 58484 32108
rect 59596 32320 59636 32360
rect 60460 36688 60500 36728
rect 60364 35932 60404 35972
rect 60172 34420 60212 34460
rect 59980 34336 60020 34376
rect 59308 32068 59348 32108
rect 58636 31816 58676 31856
rect 59116 31732 59156 31772
rect 59020 31648 59060 31688
rect 59020 31312 59060 31352
rect 58540 31060 58580 31100
rect 58348 30052 58388 30092
rect 58828 30052 58868 30092
rect 57004 29884 57044 29924
rect 56716 29800 56756 29840
rect 58828 29800 58868 29840
rect 56428 28708 56468 28748
rect 56044 28120 56084 28160
rect 55852 27868 55892 27908
rect 55180 27532 55220 27572
rect 55181 27280 55221 27320
rect 54988 26020 55028 26060
rect 55084 25936 55124 25976
rect 55372 27448 55412 27488
rect 55468 27028 55508 27068
rect 55660 27028 55700 27068
rect 55564 26608 55604 26648
rect 55756 26944 55796 26984
rect 55948 26776 55988 26816
rect 57580 29464 57620 29504
rect 57196 29380 57236 29420
rect 56908 28624 56948 28664
rect 56908 28288 56948 28328
rect 56428 27616 56468 27656
rect 56812 27532 56852 27572
rect 56332 26776 56372 26816
rect 56044 26356 56084 26396
rect 55564 26104 55604 26144
rect 54796 25852 54836 25892
rect 55660 25936 55700 25976
rect 55468 25264 55508 25304
rect 54796 24928 54836 24968
rect 54316 24508 54356 24548
rect 55276 24424 55316 24464
rect 52972 23752 53012 23792
rect 53644 23752 53684 23792
rect 54796 23752 54836 23792
rect 55756 25264 55796 25304
rect 56524 25936 56564 25976
rect 52300 22996 52340 23036
rect 52012 22828 52052 22868
rect 52108 22240 52148 22280
rect 52396 22744 52436 22784
rect 54124 23668 54164 23708
rect 52876 23416 52916 23456
rect 52972 23332 53012 23372
rect 52588 23248 52628 23288
rect 52876 23164 52916 23204
rect 52684 23080 52724 23120
rect 52780 22912 52820 22952
rect 52300 22156 52340 22196
rect 52684 22240 52724 22280
rect 52012 18460 52052 18500
rect 51436 15856 51476 15896
rect 51628 15772 51668 15812
rect 51148 15604 51188 15644
rect 51052 15520 51092 15560
rect 50572 14344 50612 14384
rect 50764 14176 50804 14216
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 51340 14176 51380 14216
rect 51244 14092 51284 14132
rect 51916 17704 51956 17744
rect 51820 15856 51860 15896
rect 51628 14344 51668 14384
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 50860 13420 50900 13460
rect 51532 13420 51572 13460
rect 50668 13168 50708 13208
rect 51628 13252 51668 13292
rect 51820 15520 51860 15560
rect 51820 13336 51860 13376
rect 51724 13084 51764 13124
rect 50380 12832 50420 12872
rect 50284 11908 50324 11948
rect 50956 12496 50996 12536
rect 52012 17284 52052 17324
rect 52012 15940 52052 15980
rect 52012 15772 52052 15812
rect 52588 21568 52628 21608
rect 54316 23164 54356 23204
rect 57004 25264 57044 25304
rect 57100 24676 57140 24716
rect 56332 24592 56372 24632
rect 55948 24508 55988 24548
rect 57388 29128 57428 29168
rect 57292 27700 57332 27740
rect 57484 25936 57524 25976
rect 57484 24508 57524 24548
rect 57196 23920 57236 23960
rect 58540 28624 58580 28664
rect 57964 28120 58004 28160
rect 58732 28120 58772 28160
rect 58060 27280 58100 27320
rect 57676 26776 57716 26816
rect 58540 27028 58580 27068
rect 58156 26944 58196 26984
rect 58348 26860 58388 26900
rect 58060 26692 58100 26732
rect 57676 26188 57716 26228
rect 57964 25768 58004 25808
rect 57676 24088 57716 24128
rect 57580 23836 57620 23876
rect 55852 23752 55892 23792
rect 56044 23752 56084 23792
rect 55276 23416 55316 23456
rect 55084 23164 55124 23204
rect 54055 22996 54095 23036
rect 53545 22912 53585 22952
rect 53655 22828 53695 22868
rect 53945 22744 53985 22784
rect 54745 22996 54785 23036
rect 54455 22744 54495 22784
rect 54855 22828 54895 22868
rect 55660 23164 55700 23204
rect 56140 23500 56180 23540
rect 56812 23752 56852 23792
rect 57292 23752 57332 23792
rect 58540 26608 58580 26648
rect 58156 25684 58196 25724
rect 58060 25096 58100 25136
rect 58060 24676 58100 24716
rect 58636 26104 58676 26144
rect 58348 25936 58388 25976
rect 58540 25936 58580 25976
rect 58444 25852 58484 25892
rect 59692 31564 59732 31604
rect 60172 33748 60212 33788
rect 60364 33244 60404 33284
rect 59788 31480 59828 31520
rect 59692 30724 59732 30764
rect 59692 30556 59732 30596
rect 59308 30052 59348 30092
rect 59404 29968 59444 30008
rect 59500 29716 59540 29756
rect 59212 29548 59252 29588
rect 59980 31648 60020 31688
rect 60076 31564 60116 31604
rect 59980 31480 60020 31520
rect 59788 30220 59828 30260
rect 59788 29800 59828 29840
rect 60076 30640 60116 30680
rect 60940 35848 60980 35888
rect 60748 32992 60788 33032
rect 60460 31732 60500 31772
rect 60460 31312 60500 31352
rect 60364 31228 60404 31268
rect 60172 29716 60212 29756
rect 60076 29632 60116 29672
rect 60268 29548 60308 29588
rect 60556 30136 60596 30176
rect 61036 34336 61076 34376
rect 63532 37948 63572 37988
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 62956 37360 62996 37400
rect 61612 37276 61652 37316
rect 61516 36940 61556 36980
rect 61420 36688 61460 36728
rect 63436 37276 63476 37316
rect 61420 36016 61460 36056
rect 62092 36520 62132 36560
rect 61228 35848 61268 35888
rect 61516 35932 61556 35972
rect 61420 35512 61460 35552
rect 61420 35008 61460 35048
rect 61324 33580 61364 33620
rect 61132 33496 61172 33536
rect 61324 32992 61364 33032
rect 61132 31816 61172 31856
rect 60748 30556 60788 30596
rect 60940 30388 60980 30428
rect 60940 30220 60980 30260
rect 60460 29464 60500 29504
rect 60652 29128 60692 29168
rect 60556 29044 60596 29084
rect 59308 28456 59348 28496
rect 58924 28036 58964 28076
rect 58828 27280 58868 27320
rect 59116 28288 59156 28328
rect 59020 27112 59060 27152
rect 58828 26944 58868 26984
rect 59020 26776 59060 26816
rect 59212 26944 59252 26984
rect 58828 26608 58868 26648
rect 59692 28288 59732 28328
rect 59596 27784 59636 27824
rect 59884 28120 59924 28160
rect 60844 29464 60884 29504
rect 61132 30640 61172 30680
rect 61132 30136 61172 30176
rect 61036 29212 61076 29252
rect 60940 29044 60980 29084
rect 60844 28540 60884 28580
rect 60172 28288 60212 28328
rect 60364 28288 60404 28328
rect 59788 28036 59828 28076
rect 60076 27868 60116 27908
rect 59884 27784 59924 27824
rect 59980 27700 60020 27740
rect 60460 28036 60500 28076
rect 60364 27868 60404 27908
rect 60748 28288 60788 28328
rect 61612 35848 61652 35888
rect 62188 36016 62228 36056
rect 62092 35848 62132 35888
rect 62668 35848 62708 35888
rect 61996 35764 62036 35804
rect 61708 35512 61748 35552
rect 61516 34672 61556 34712
rect 62188 34756 62228 34796
rect 61900 34504 61940 34544
rect 62092 34336 62132 34376
rect 62092 34000 62132 34040
rect 61612 33664 61652 33704
rect 61516 32992 61556 33032
rect 61612 32068 61652 32108
rect 61900 32068 61940 32108
rect 61900 31648 61940 31688
rect 61420 29884 61460 29924
rect 61324 29632 61364 29672
rect 61228 29128 61268 29168
rect 61612 29464 61652 29504
rect 61516 28540 61556 28580
rect 62668 34756 62708 34796
rect 63532 37192 63572 37232
rect 63532 36688 63572 36728
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 62572 34504 62612 34544
rect 62668 34420 62708 34460
rect 62764 34336 62804 34376
rect 62668 34252 62708 34292
rect 62572 34000 62612 34040
rect 62380 33664 62420 33704
rect 62860 34000 62900 34040
rect 62188 33580 62228 33620
rect 62092 31312 62132 31352
rect 62476 33496 62516 33536
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 63244 34420 63284 34460
rect 63052 34252 63092 34292
rect 70156 38284 70196 38324
rect 71404 38284 71444 38324
rect 63820 36688 63860 36728
rect 63724 36520 63764 36560
rect 67468 38200 67508 38240
rect 64300 37948 64340 37988
rect 65548 37360 65588 37400
rect 64204 37276 64244 37316
rect 64108 37192 64148 37232
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 64012 36688 64052 36728
rect 63628 34420 63668 34460
rect 63244 34084 63284 34124
rect 63148 34000 63188 34040
rect 63052 33748 63092 33788
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 62476 32908 62516 32948
rect 62284 32824 62324 32864
rect 62572 32824 62612 32864
rect 62860 33076 62900 33116
rect 62476 32068 62516 32108
rect 62668 32488 62708 32528
rect 64108 36520 64148 36560
rect 65548 36688 65588 36728
rect 66316 37360 66356 37400
rect 65740 36436 65780 36476
rect 64204 35764 64244 35804
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 66028 35680 66068 35720
rect 65164 35596 65204 35636
rect 64108 34672 64148 34712
rect 63052 32236 63092 32276
rect 64108 33076 64148 33116
rect 64012 32908 64052 32948
rect 63436 32488 63476 32528
rect 63244 32236 63284 32276
rect 62860 31900 62900 31940
rect 63532 31900 63572 31940
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 65836 35344 65876 35384
rect 65932 35008 65972 35048
rect 65452 34084 65492 34124
rect 65932 33496 65972 33536
rect 66124 35176 66164 35216
rect 66700 37276 66740 37316
rect 66988 36688 67028 36728
rect 67276 37360 67316 37400
rect 67084 36184 67124 36224
rect 66700 35932 66740 35972
rect 66988 35848 67028 35888
rect 67372 36856 67412 36896
rect 67756 38032 67796 38072
rect 67756 37612 67796 37652
rect 68236 37612 68276 37652
rect 67948 37276 67988 37316
rect 67564 37108 67604 37148
rect 67756 36520 67796 36560
rect 67564 36268 67604 36308
rect 66892 35764 66932 35804
rect 66796 35344 66836 35384
rect 66892 35260 66932 35300
rect 66604 35176 66644 35216
rect 66412 34504 66452 34544
rect 66220 34168 66260 34208
rect 66796 35176 66836 35216
rect 66700 34588 66740 34628
rect 66316 33916 66356 33956
rect 66700 34420 66740 34460
rect 66124 33580 66164 33620
rect 66220 33496 66260 33536
rect 64108 32236 64148 32276
rect 64012 31900 64052 31940
rect 62668 31228 62708 31268
rect 63052 31312 63092 31352
rect 63358 31396 63398 31436
rect 62476 30640 62516 30680
rect 62284 30556 62324 30596
rect 62860 30640 62900 30680
rect 61708 29212 61748 29252
rect 63724 30640 63764 30680
rect 63820 30556 63860 30596
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 63244 30052 63284 30092
rect 63340 29968 63380 30008
rect 63436 29800 63476 29840
rect 63052 29632 63092 29672
rect 63532 29548 63572 29588
rect 63436 29296 63476 29336
rect 63052 29212 63092 29252
rect 63916 29800 63956 29840
rect 60844 28036 60884 28076
rect 58924 26104 58964 26144
rect 59404 26104 59444 26144
rect 59308 26020 59348 26060
rect 59212 25936 59252 25976
rect 58828 25768 58868 25808
rect 58636 24844 58676 24884
rect 59020 25684 59060 25724
rect 59020 25516 59060 25556
rect 58828 25096 58868 25136
rect 58732 24676 58772 24716
rect 58924 24844 58964 24884
rect 56428 23248 56468 23288
rect 56455 22996 56495 23036
rect 56812 23248 56852 23288
rect 57292 23416 57332 23456
rect 57676 23584 57716 23624
rect 58060 23584 58100 23624
rect 57655 22744 57695 22784
rect 60172 27448 60212 27488
rect 60652 27448 60692 27488
rect 60076 27364 60116 27404
rect 59788 26524 59828 26564
rect 59596 25264 59636 25304
rect 59404 25096 59444 25136
rect 59596 24844 59636 24884
rect 60460 27196 60500 27236
rect 60364 26860 60404 26900
rect 60268 26776 60308 26816
rect 59788 25936 59828 25976
rect 60172 25600 60212 25640
rect 59884 25096 59924 25136
rect 59788 24844 59828 24884
rect 60172 24844 60212 24884
rect 59500 24760 59540 24800
rect 59404 24676 59444 24716
rect 60076 24760 60116 24800
rect 60748 27112 60788 27152
rect 61228 28372 61268 28412
rect 61420 27952 61460 27992
rect 61132 27196 61172 27236
rect 61036 27112 61076 27152
rect 60748 26860 60788 26900
rect 60556 26692 60596 26732
rect 61324 26608 61364 26648
rect 60940 26524 60980 26564
rect 60556 26440 60596 26480
rect 60364 26188 60404 26228
rect 61132 26440 61172 26480
rect 61132 26188 61172 26228
rect 60460 26104 60500 26144
rect 60556 26020 60596 26060
rect 60748 26020 60788 26060
rect 60364 25852 60404 25892
rect 60748 25768 60788 25808
rect 60940 25348 60980 25388
rect 60460 25096 60500 25136
rect 60844 23920 60884 23960
rect 61228 23920 61268 23960
rect 60460 23836 60500 23876
rect 60748 23836 60788 23876
rect 58444 23164 58484 23204
rect 59020 23752 59060 23792
rect 58828 23164 58868 23204
rect 59692 23752 59732 23792
rect 59980 23752 60020 23792
rect 59308 23500 59348 23540
rect 59692 23500 59732 23540
rect 59020 22744 59060 22784
rect 59255 22744 59295 22784
rect 60076 23584 60116 23624
rect 61420 26104 61460 26144
rect 61612 28372 61652 28412
rect 61804 28288 61844 28328
rect 61900 27784 61940 27824
rect 61612 26608 61652 26648
rect 61612 26440 61652 26480
rect 61612 26188 61652 26228
rect 61900 27028 61940 27068
rect 61900 26776 61940 26816
rect 61804 26104 61844 26144
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 63148 28288 63188 28328
rect 64012 29296 64052 29336
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 64492 32320 64532 32360
rect 64780 32236 64820 32276
rect 64300 31984 64340 32024
rect 64204 31648 64244 31688
rect 64396 31396 64436 31436
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 65164 31900 65204 31940
rect 64396 30640 64436 30680
rect 64204 30556 64244 30596
rect 64780 29800 64820 29840
rect 64204 29464 64244 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 63820 28204 63860 28244
rect 64012 29128 64052 29168
rect 62860 26776 62900 26816
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 63916 27784 63956 27824
rect 63820 27616 63860 27656
rect 64204 29128 64244 29168
rect 64780 29128 64820 29168
rect 65068 28792 65108 28832
rect 64300 28204 64340 28244
rect 64780 28288 64820 28328
rect 65164 28456 65204 28496
rect 66028 32824 66068 32864
rect 66796 34168 66836 34208
rect 65644 32656 65684 32696
rect 65356 32488 65396 32528
rect 65932 32572 65972 32612
rect 65644 32320 65684 32360
rect 65356 32236 65396 32276
rect 65452 31984 65492 32024
rect 66220 32404 66260 32444
rect 66124 31900 66164 31940
rect 65836 30724 65876 30764
rect 65356 30220 65396 30260
rect 65548 30220 65588 30260
rect 65932 30556 65972 30596
rect 66124 30724 66164 30764
rect 65452 29800 65492 29840
rect 65836 29800 65876 29840
rect 65644 29296 65684 29336
rect 65548 28792 65588 28832
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 65260 28120 65300 28160
rect 65068 28036 65108 28076
rect 64876 27784 64916 27824
rect 64876 27616 64916 27656
rect 63628 26944 63668 26984
rect 64204 26944 64244 26984
rect 64012 26860 64052 26900
rect 63820 26776 63860 26816
rect 62956 26524 62996 26564
rect 63532 26272 63572 26312
rect 62860 26104 62900 26144
rect 61516 25852 61556 25892
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 64012 26524 64052 26564
rect 63820 26104 63860 26144
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 64396 26272 64436 26312
rect 65164 27952 65204 27992
rect 65356 27616 65396 27656
rect 65452 27532 65492 27572
rect 65260 27364 65300 27404
rect 65164 27280 65204 27320
rect 64780 26188 64820 26228
rect 64300 25936 64340 25976
rect 64780 25936 64820 25976
rect 64972 25936 65012 25976
rect 63148 25264 63188 25304
rect 61516 25096 61556 25136
rect 61708 25012 61748 25052
rect 62572 24760 62612 24800
rect 62476 24256 62516 24296
rect 62092 24004 62132 24044
rect 62572 24004 62612 24044
rect 63436 25264 63476 25304
rect 63532 25096 63572 25136
rect 63436 24928 63476 24968
rect 63244 23920 63284 23960
rect 63628 24592 63668 24632
rect 63916 25264 63956 25304
rect 63916 24844 63956 24884
rect 65068 25684 65108 25724
rect 63916 24676 63956 24716
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 64108 24592 64148 24632
rect 64588 24676 64628 24716
rect 64396 24592 64436 24632
rect 64492 24424 64532 24464
rect 65068 25096 65108 25136
rect 65836 29128 65876 29168
rect 65740 28036 65780 28076
rect 67372 35848 67412 35888
rect 67276 35260 67316 35300
rect 66988 34672 67028 34712
rect 67468 34672 67508 34712
rect 67660 34588 67700 34628
rect 66892 32488 66932 32528
rect 66892 32320 66932 32360
rect 66604 31984 66644 32024
rect 66412 31396 66452 31436
rect 66796 31396 66836 31436
rect 66700 31228 66740 31268
rect 66604 31060 66644 31100
rect 66316 28792 66356 28832
rect 65644 27952 65684 27992
rect 65932 27952 65972 27992
rect 65836 27616 65876 27656
rect 65740 27532 65780 27572
rect 65548 26524 65588 26564
rect 65356 26104 65396 26144
rect 65356 25936 65396 25976
rect 62476 23584 62516 23624
rect 65644 26104 65684 26144
rect 65548 24592 65588 24632
rect 65260 23920 65300 23960
rect 65644 23920 65684 23960
rect 63244 23668 63284 23708
rect 63628 23668 63668 23708
rect 62860 23584 62900 23624
rect 62764 23332 62804 23372
rect 60464 22744 60504 22784
rect 63244 23332 63284 23372
rect 64108 23752 64148 23792
rect 65932 26524 65972 26564
rect 66124 27952 66164 27992
rect 66028 23920 66068 23960
rect 66412 26776 66452 26816
rect 66316 25348 66356 25388
rect 66412 24928 66452 24968
rect 66412 24676 66452 24716
rect 67276 34336 67316 34376
rect 67180 34168 67220 34208
rect 67180 33916 67220 33956
rect 67180 32320 67220 32360
rect 67084 31900 67124 31940
rect 66988 31396 67028 31436
rect 66988 31228 67028 31268
rect 67084 31060 67124 31100
rect 67276 30640 67316 30680
rect 66796 29296 66836 29336
rect 66892 28624 66932 28664
rect 66796 28288 66836 28328
rect 66796 27364 66836 27404
rect 66796 25264 66836 25304
rect 66700 25012 66740 25052
rect 66700 24676 66740 24716
rect 67564 34336 67604 34376
rect 67669 34336 67709 34376
rect 67468 34252 67508 34292
rect 68140 37276 68180 37316
rect 68140 36856 68180 36896
rect 68044 35512 68084 35552
rect 68428 37276 68468 37316
rect 68332 37192 68372 37232
rect 68716 37780 68756 37820
rect 69388 38116 69428 38156
rect 69388 37780 69428 37820
rect 68716 36688 68756 36728
rect 69196 36940 69236 36980
rect 69100 36856 69140 36896
rect 68716 36520 68756 36560
rect 68428 36436 68468 36476
rect 69004 36436 69044 36476
rect 68716 36016 68756 36056
rect 68524 35932 68564 35972
rect 68236 35176 68276 35216
rect 68044 34504 68084 34544
rect 67564 33916 67604 33956
rect 67468 28960 67508 29000
rect 66988 28288 67028 28328
rect 67372 28288 67412 28328
rect 67852 31816 67892 31856
rect 67660 29632 67700 29672
rect 67564 27532 67604 27572
rect 67276 26440 67316 26480
rect 67180 26104 67220 26144
rect 67660 26776 67700 26816
rect 67756 26524 67796 26564
rect 67948 30640 67988 30680
rect 68332 29800 68372 29840
rect 68236 29716 68276 29756
rect 68044 28960 68084 29000
rect 68428 29212 68468 29252
rect 68332 28792 68372 28832
rect 68140 28036 68180 28076
rect 68140 27616 68180 27656
rect 68332 27448 68372 27488
rect 68812 35680 68852 35720
rect 68908 34588 68948 34628
rect 69292 36856 69332 36896
rect 69484 37192 69524 37232
rect 69484 36772 69524 36812
rect 70540 36856 70580 36896
rect 69772 36688 69812 36728
rect 69100 36352 69140 36392
rect 69100 36184 69140 36224
rect 69004 34420 69044 34460
rect 68620 32824 68660 32864
rect 68620 31480 68660 31520
rect 68812 32824 68852 32864
rect 69196 34840 69236 34880
rect 69004 32656 69044 32696
rect 69100 32488 69140 32528
rect 68908 32404 68948 32444
rect 68812 31480 68852 31520
rect 68908 30640 68948 30680
rect 68524 27364 68564 27404
rect 68428 26776 68468 26816
rect 68044 26524 68084 26564
rect 68428 26356 68468 26396
rect 67852 26272 67892 26312
rect 67372 26188 67412 26228
rect 67084 25348 67124 25388
rect 67852 25852 67892 25892
rect 68236 25852 68276 25892
rect 68140 25684 68180 25724
rect 68620 26104 68660 26144
rect 67660 25012 67700 25052
rect 67372 24760 67412 24800
rect 67852 25012 67892 25052
rect 67660 24676 67700 24716
rect 68332 24760 68372 24800
rect 68140 24592 68180 24632
rect 67276 24508 67316 24548
rect 67756 24004 67796 24044
rect 67276 23752 67316 23792
rect 67660 23752 67700 23792
rect 68524 23920 68564 23960
rect 69100 31060 69140 31100
rect 69100 29800 69140 29840
rect 68908 27868 68948 27908
rect 69292 32320 69332 32360
rect 69292 29968 69332 30008
rect 69676 36184 69716 36224
rect 69484 36100 69524 36140
rect 70060 36520 70100 36560
rect 70060 36016 70100 36056
rect 69868 35848 69908 35888
rect 69964 34588 70004 34628
rect 69868 34336 69908 34376
rect 71116 37192 71156 37232
rect 71500 37192 71540 37232
rect 71980 37024 72020 37064
rect 71116 36772 71156 36812
rect 70636 36520 70676 36560
rect 70924 36436 70964 36476
rect 70924 36100 70964 36140
rect 70540 35428 70580 35468
rect 70828 35428 70868 35468
rect 70444 35260 70484 35300
rect 70540 35176 70580 35216
rect 70444 34588 70484 34628
rect 70348 34504 70388 34544
rect 69580 34084 69620 34124
rect 69484 31648 69524 31688
rect 69484 30640 69524 30680
rect 69484 30052 69524 30092
rect 69484 27868 69524 27908
rect 69868 33916 69908 33956
rect 70348 33160 70388 33200
rect 69772 32656 69812 32696
rect 69676 32488 69716 32528
rect 69964 32320 70004 32360
rect 70732 35176 70772 35216
rect 70636 34504 70676 34544
rect 71020 35512 71060 35552
rect 69868 31984 69908 32024
rect 70540 32656 70580 32696
rect 70636 31648 70676 31688
rect 70828 32656 70868 32696
rect 70924 32404 70964 32444
rect 72076 36520 72116 36560
rect 72172 36436 72212 36476
rect 71212 36100 71252 36140
rect 71884 36100 71924 36140
rect 71116 32908 71156 32948
rect 71116 32488 71156 32528
rect 71020 32320 71060 32360
rect 71116 32236 71156 32276
rect 70732 31564 70772 31604
rect 70444 31144 70484 31184
rect 70924 31396 70964 31436
rect 70732 31312 70772 31352
rect 70828 31144 70868 31184
rect 69772 29548 69812 29588
rect 69964 29632 70004 29672
rect 70636 30724 70676 30764
rect 70540 30640 70580 30680
rect 70540 30052 70580 30092
rect 70540 29800 70580 29840
rect 70732 30052 70772 30092
rect 70252 29548 70292 29588
rect 70060 29464 70100 29504
rect 70636 29464 70676 29504
rect 70444 29128 70484 29168
rect 70060 29044 70100 29084
rect 70540 29044 70580 29084
rect 70252 28960 70292 29000
rect 71116 31564 71156 31604
rect 71116 31144 71156 31184
rect 71596 35848 71636 35888
rect 72556 36352 72596 36392
rect 71980 35848 72020 35888
rect 71404 35260 71444 35300
rect 71308 34504 71348 34544
rect 71404 34168 71444 34208
rect 71884 35176 71924 35216
rect 71692 35008 71732 35048
rect 72556 35260 72596 35300
rect 72364 35008 72404 35048
rect 72556 35008 72596 35048
rect 72076 34924 72116 34964
rect 72460 34924 72500 34964
rect 71788 34504 71828 34544
rect 71980 34336 72020 34376
rect 71788 34168 71828 34208
rect 71596 33664 71636 33704
rect 73036 37444 73076 37484
rect 72940 37192 72980 37232
rect 72940 37024 72980 37064
rect 72844 36688 72884 36728
rect 72748 36436 72788 36476
rect 72748 35176 72788 35216
rect 72748 35008 72788 35048
rect 71980 33832 72020 33872
rect 71692 32656 71732 32696
rect 71500 32404 71540 32444
rect 71596 32320 71636 32360
rect 71308 31312 71348 31352
rect 70924 30136 70964 30176
rect 71020 29800 71060 29840
rect 71212 30808 71252 30848
rect 71308 30724 71348 30764
rect 71404 30472 71444 30512
rect 71212 30388 71252 30428
rect 72460 33664 72500 33704
rect 72268 33580 72308 33620
rect 72556 33580 72596 33620
rect 72556 32824 72596 32864
rect 71980 32656 72020 32696
rect 71884 32320 71924 32360
rect 72076 32488 72116 32528
rect 71692 30220 71732 30260
rect 70924 29716 70964 29756
rect 70924 29380 70964 29420
rect 70732 29128 70772 29168
rect 71116 29044 71156 29084
rect 72652 32320 72692 32360
rect 72940 36436 72980 36476
rect 73036 35932 73076 35972
rect 73612 37444 73652 37484
rect 73228 37360 73268 37400
rect 73420 37276 73460 37316
rect 73996 37360 74036 37400
rect 73900 37276 73940 37316
rect 73228 36856 73268 36896
rect 73324 36772 73364 36812
rect 73516 36520 73556 36560
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 73804 36772 73844 36812
rect 74092 36940 74132 36980
rect 74380 37276 74420 37316
rect 74764 37360 74804 37400
rect 74572 37192 74612 37232
rect 75052 37192 75092 37232
rect 76780 37360 76820 37400
rect 75244 36856 75284 36896
rect 74476 36184 74516 36224
rect 74284 36100 74324 36140
rect 75148 36688 75188 36728
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 76588 36772 76628 36812
rect 76204 36688 76244 36728
rect 75244 36520 75284 36560
rect 76108 36520 76148 36560
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 73516 36016 73556 36056
rect 73036 35260 73076 35300
rect 72844 32824 72884 32864
rect 72172 31984 72212 32024
rect 72748 32152 72788 32192
rect 72652 32068 72692 32108
rect 72556 31984 72596 32024
rect 72364 31732 72404 31772
rect 72172 30388 72212 30428
rect 72076 30136 72116 30176
rect 71404 29800 71444 29840
rect 71308 29716 71348 29756
rect 71788 29800 71828 29840
rect 71980 29884 72020 29924
rect 72076 29800 72116 29840
rect 72268 30136 72308 30176
rect 72268 29380 72308 29420
rect 71884 29296 71924 29336
rect 71308 28960 71348 29000
rect 70828 28876 70868 28916
rect 71212 28876 71252 28916
rect 69388 27784 69428 27824
rect 68908 27448 68948 27488
rect 68812 27196 68852 27236
rect 69004 27196 69044 27236
rect 68908 26776 68948 26816
rect 68812 26524 68852 26564
rect 69004 26272 69044 26312
rect 68908 23920 68948 23960
rect 68716 23752 68756 23792
rect 70060 27700 70100 27740
rect 69388 26440 69428 26480
rect 69292 26104 69332 26144
rect 69772 27616 69812 27656
rect 69772 27448 69812 27488
rect 69484 26188 69524 26228
rect 69196 25264 69236 25304
rect 70252 27700 70292 27740
rect 70540 28288 70580 28328
rect 70636 28120 70676 28160
rect 70540 27868 70580 27908
rect 70252 27364 70292 27404
rect 70444 26608 70484 26648
rect 72940 32488 72980 32528
rect 72940 32320 72980 32360
rect 73228 35092 73268 35132
rect 73132 32908 73172 32948
rect 73036 32068 73076 32108
rect 72940 31816 72980 31856
rect 73036 31648 73076 31688
rect 73036 31312 73076 31352
rect 72652 30472 72692 30512
rect 72460 30220 72500 30260
rect 72556 29380 72596 29420
rect 71500 29128 71540 29168
rect 72460 29128 72500 29168
rect 70828 28120 70868 28160
rect 71980 29044 72020 29084
rect 71884 28876 71924 28916
rect 71692 28372 71732 28412
rect 71500 27868 71540 27908
rect 71500 27700 71540 27740
rect 71308 27364 71348 27404
rect 70828 27280 70868 27320
rect 71404 27280 71444 27320
rect 70348 25264 70388 25304
rect 70348 25096 70388 25136
rect 70924 26608 70964 26648
rect 71308 26272 71348 26312
rect 70540 24844 70580 24884
rect 70348 24760 70388 24800
rect 71308 26104 71348 26144
rect 71212 25432 71252 25472
rect 71020 24592 71060 24632
rect 70156 23920 70196 23960
rect 70540 23920 70580 23960
rect 70828 23920 70868 23960
rect 68908 23584 68948 23624
rect 69292 23584 69332 23624
rect 70156 23752 70196 23792
rect 70444 23752 70484 23792
rect 71788 27616 71828 27656
rect 71596 27364 71636 27404
rect 71596 26272 71636 26312
rect 71788 26272 71828 26312
rect 72364 26692 72404 26732
rect 71980 26608 72020 26648
rect 72556 26440 72596 26480
rect 72556 26188 72596 26228
rect 71980 26104 72020 26144
rect 73036 26860 73076 26900
rect 72652 25852 72692 25892
rect 71788 25432 71828 25472
rect 71596 24760 71636 24800
rect 71692 24592 71732 24632
rect 72844 25432 72884 25472
rect 73036 25432 73076 25472
rect 71884 25264 71924 25304
rect 72652 25264 72692 25304
rect 72460 25096 72500 25136
rect 72076 24928 72116 24968
rect 70924 23752 70964 23792
rect 71692 23752 71732 23792
rect 71980 23752 72020 23792
rect 73420 35848 73460 35888
rect 73804 35932 73844 35972
rect 73996 35848 74036 35888
rect 74284 35596 74324 35636
rect 73708 35428 73748 35468
rect 74188 35176 74228 35216
rect 73708 33916 73748 33956
rect 73324 31648 73364 31688
rect 73516 31060 73556 31100
rect 73228 29044 73268 29084
rect 73420 28540 73460 28580
rect 73612 30808 73652 30848
rect 73708 30388 73748 30428
rect 73516 27616 73556 27656
rect 73228 25936 73268 25976
rect 73132 24172 73172 24212
rect 73324 23920 73364 23960
rect 73612 23920 73652 23960
rect 74764 36016 74804 36056
rect 75436 36016 75476 36056
rect 75916 35932 75956 35972
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 74572 34168 74612 34208
rect 75628 34168 75668 34208
rect 74860 33664 74900 33704
rect 74764 33412 74804 33452
rect 74860 33160 74900 33200
rect 74572 31816 74612 31856
rect 75532 33496 75572 33536
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 74284 31732 74324 31772
rect 74188 30388 74228 30428
rect 73804 28372 73844 28412
rect 73900 27616 73940 27656
rect 73900 24004 73940 24044
rect 74092 27364 74132 27404
rect 74284 26104 74324 26144
rect 74476 26272 74516 26312
rect 74476 25936 74516 25976
rect 74380 25852 74420 25892
rect 74860 31648 74900 31688
rect 74668 31312 74708 31352
rect 74860 30724 74900 30764
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 75436 30808 75476 30848
rect 75820 33580 75860 33620
rect 76300 36604 76340 36644
rect 76876 36688 76916 36728
rect 76780 36604 76820 36644
rect 76588 36520 76628 36560
rect 76684 36184 76724 36224
rect 76492 35848 76532 35888
rect 76780 36100 76820 36140
rect 77164 37360 77204 37400
rect 77452 37360 77492 37400
rect 77260 37192 77300 37232
rect 77356 36772 77396 36812
rect 77068 36520 77108 36560
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 76108 35176 76148 35216
rect 76492 35008 76532 35048
rect 77068 35596 77108 35636
rect 77164 35344 77204 35384
rect 76876 35008 76916 35048
rect 76204 34336 76244 34376
rect 77548 36100 77588 36140
rect 77932 37192 77972 37232
rect 77452 35596 77492 35636
rect 77644 35344 77684 35384
rect 77452 35176 77492 35216
rect 78508 37360 78548 37400
rect 78316 37276 78356 37316
rect 79468 37276 79508 37316
rect 78220 36688 78260 36728
rect 78316 36016 78356 36056
rect 78124 35428 78164 35468
rect 77836 35176 77876 35216
rect 78124 34588 78164 34628
rect 77644 34336 77684 34376
rect 77932 34336 77972 34376
rect 78124 34336 78164 34376
rect 79468 34336 79508 34376
rect 76876 34252 76916 34292
rect 77356 34252 77396 34292
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 77260 33832 77300 33872
rect 76876 33748 76916 33788
rect 76300 33664 76340 33704
rect 76492 33664 76532 33704
rect 76396 33496 76436 33536
rect 76012 33412 76052 33452
rect 76012 32320 76052 32360
rect 75820 32152 75860 32192
rect 75340 30724 75380 30764
rect 75148 30640 75188 30680
rect 75532 30556 75572 30596
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 75052 29884 75092 29924
rect 75436 30052 75476 30092
rect 75820 30052 75860 30092
rect 76012 32152 76052 32192
rect 76972 33664 77012 33704
rect 76780 33412 76820 33452
rect 76588 32656 76628 32696
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 76300 32320 76340 32360
rect 76492 32320 76532 32360
rect 76204 31648 76244 31688
rect 76204 31480 76244 31520
rect 76108 31144 76148 31184
rect 76684 32236 76724 32276
rect 77164 32824 77204 32864
rect 76876 32152 76916 32192
rect 76492 31480 76532 31520
rect 77452 33664 77492 33704
rect 78412 33664 78452 33704
rect 77548 33412 77588 33452
rect 77452 32320 77492 32360
rect 77836 32824 77876 32864
rect 78124 32824 78164 32864
rect 78508 32824 78548 32864
rect 77740 32152 77780 32192
rect 76780 31312 76820 31352
rect 76012 30640 76052 30680
rect 76300 31144 76340 31184
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 76492 30724 76532 30764
rect 76108 30220 76148 30260
rect 75628 29884 75668 29924
rect 75532 29800 75572 29840
rect 74860 29632 74900 29672
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 75340 28540 75380 28580
rect 75436 28288 75476 28328
rect 75244 27700 75284 27740
rect 75052 27616 75092 27656
rect 75244 27364 75284 27404
rect 75820 29716 75860 29756
rect 76012 29800 76052 29840
rect 75916 29632 75956 29672
rect 75820 29212 75860 29252
rect 76588 30640 76628 30680
rect 76492 30472 76532 30512
rect 76780 30472 76820 30512
rect 77164 31312 77204 31352
rect 77068 31228 77108 31268
rect 77452 31144 77492 31184
rect 77164 31060 77204 31100
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 76684 29296 76724 29336
rect 76492 29212 76532 29252
rect 76108 28960 76148 29000
rect 76396 28372 76436 28412
rect 76780 28624 76820 28664
rect 77452 30640 77492 30680
rect 77644 30724 77684 30764
rect 77644 30472 77684 30512
rect 77260 30220 77300 30260
rect 77260 29632 77300 29672
rect 77068 29296 77108 29336
rect 77068 28624 77108 28664
rect 76876 28288 76916 28328
rect 77452 28288 77492 28328
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 75436 27700 75476 27740
rect 74860 26860 74900 26900
rect 74764 26776 74804 26816
rect 74764 26356 74804 26396
rect 74668 26272 74708 26312
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 75148 27028 75188 27068
rect 75340 27028 75380 27068
rect 74860 26188 74900 26228
rect 74860 25936 74900 25976
rect 75436 26860 75476 26900
rect 75436 25936 75476 25976
rect 74476 25264 74516 25304
rect 74572 25180 74612 25220
rect 74476 24760 74516 24800
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 75436 25348 75476 25388
rect 74956 24760 74996 24800
rect 73804 23920 73844 23960
rect 73996 23920 74036 23960
rect 75244 24172 75284 24212
rect 74476 24004 74516 24044
rect 74860 23920 74900 23960
rect 74476 23248 74516 23288
rect 75628 27028 75668 27068
rect 75724 26944 75764 26984
rect 75628 26776 75668 26816
rect 75628 26524 75668 26564
rect 75724 26356 75764 26396
rect 75916 26776 75956 26816
rect 76588 26776 76628 26816
rect 76204 26608 76244 26648
rect 76492 26608 76532 26648
rect 76780 27616 76820 27656
rect 76972 27616 77012 27656
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 76876 26272 76916 26312
rect 75628 25936 75668 25976
rect 75820 26188 75860 26228
rect 75916 26104 75956 26144
rect 76396 26104 76436 26144
rect 75820 25936 75860 25976
rect 75724 25348 75764 25388
rect 76204 25852 76244 25892
rect 75724 24592 75764 24632
rect 76684 25936 76724 25976
rect 77164 27448 77204 27488
rect 77068 26272 77108 26312
rect 77356 26608 77396 26648
rect 79468 32152 79508 32192
rect 78316 31648 78356 31688
rect 78220 31312 78260 31352
rect 77836 30640 77876 30680
rect 77836 30472 77876 30512
rect 79468 30472 79508 30512
rect 77836 28708 77876 28748
rect 78124 28288 78164 28328
rect 79468 28288 79508 28328
rect 76780 25852 76820 25892
rect 76300 25180 76340 25220
rect 76684 25180 76724 25220
rect 76204 24928 76244 24968
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 76492 24760 76532 24800
rect 76684 24592 76724 24632
rect 76108 23752 76148 23792
rect 76492 23752 76532 23792
rect 76972 23752 77012 23792
rect 77836 25852 77876 25892
rect 74860 23416 74900 23456
rect 74860 23248 74900 23288
rect 75244 23584 75284 23624
rect 75244 23416 75284 23456
rect 75628 23584 75668 23624
rect 77932 25264 77972 25304
rect 78508 26608 78548 26648
rect 79468 26608 79508 26648
rect 78316 25264 78356 25304
rect 78988 24592 79028 24632
rect 77452 23752 77492 23792
rect 79084 23752 79124 23792
rect 78796 23416 78836 23456
rect 79276 23416 79316 23456
rect 78604 22744 78644 22784
rect 78855 22744 78895 22784
rect 52972 21988 53012 22028
rect 52588 20140 52628 20180
rect 52300 18544 52340 18584
rect 52396 17284 52436 17324
rect 52780 18124 52820 18164
rect 52684 17200 52724 17240
rect 52300 17116 52340 17156
rect 52492 17116 52532 17156
rect 52204 17032 52244 17072
rect 52396 16948 52436 16988
rect 52588 17032 52628 17072
rect 52204 16780 52244 16820
rect 53836 17200 53876 17240
rect 53655 17116 53695 17156
rect 54437 17284 54477 17324
rect 54345 17200 54385 17240
rect 54055 17116 54095 17156
rect 54508 17116 54548 17156
rect 53932 17032 53972 17072
rect 54412 17032 54452 17072
rect 53836 16528 53876 16568
rect 52780 16192 52820 16232
rect 52108 14428 52148 14468
rect 52588 15520 52628 15560
rect 52492 15268 52532 15308
rect 52300 14680 52340 14720
rect 52972 15856 53012 15896
rect 53164 15856 53204 15896
rect 52780 15688 52820 15728
rect 53452 15856 53492 15896
rect 53164 15688 53204 15728
rect 52684 14512 52724 14552
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 52204 14176 52244 14216
rect 52972 14092 53012 14132
rect 53164 15436 53204 15476
rect 53356 15268 53396 15308
rect 54855 17200 54895 17240
rect 55145 17200 55185 17240
rect 54745 17032 54785 17072
rect 55468 16696 55508 16736
rect 54796 16192 54836 16232
rect 55660 16612 55700 16652
rect 55948 16612 55988 16652
rect 56524 16192 56564 16232
rect 56140 16024 56180 16064
rect 55468 15940 55508 15980
rect 54604 15772 54644 15812
rect 53644 15604 53684 15644
rect 53068 13840 53108 13880
rect 53836 14008 53876 14048
rect 54412 14428 54452 14468
rect 53548 13588 53588 13628
rect 53452 13420 53492 13460
rect 53260 13168 53300 13208
rect 54508 13672 54548 13712
rect 51916 12832 51956 12872
rect 51820 12664 51860 12704
rect 51820 12496 51860 12536
rect 50764 11908 50804 11948
rect 50380 11740 50420 11780
rect 50188 11572 50228 11612
rect 49996 10984 50036 11024
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 51148 11572 51188 11612
rect 50380 11488 50420 11528
rect 50860 11068 50900 11108
rect 51340 10984 51380 11024
rect 51820 12076 51860 12116
rect 52012 12076 52052 12116
rect 51916 11656 51956 11696
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 52204 11824 52244 11864
rect 52108 11656 52148 11696
rect 52108 11488 52148 11528
rect 50668 10648 50708 10688
rect 50284 10312 50324 10352
rect 49900 9640 49940 9680
rect 49900 9136 49940 9176
rect 49228 8800 49268 8840
rect 49132 8632 49172 8672
rect 49036 8548 49076 8588
rect 48844 8296 48884 8336
rect 48940 8128 48980 8168
rect 48844 7999 48884 8000
rect 48844 7960 48884 7999
rect 49228 7960 49268 8000
rect 48748 7792 48788 7832
rect 48364 7372 48404 7412
rect 48556 5860 48596 5900
rect 48460 5692 48500 5732
rect 48364 5524 48404 5564
rect 47884 5440 47924 5480
rect 48268 4936 48308 4976
rect 48556 5020 48596 5060
rect 48460 4936 48500 4976
rect 49036 7624 49076 7664
rect 48748 5860 48788 5900
rect 49804 8632 49844 8672
rect 50764 9136 50804 9176
rect 49996 8632 50036 8672
rect 50188 8548 50228 8588
rect 49900 8212 49940 8252
rect 49708 7708 49748 7748
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 51532 8800 51572 8840
rect 51340 8632 51380 8672
rect 51628 8716 51668 8756
rect 52012 10312 52052 10352
rect 51916 8884 51956 8924
rect 51820 8800 51860 8840
rect 51724 8464 51764 8504
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 50476 7204 50516 7244
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 52300 9976 52340 10016
rect 52108 9556 52148 9596
rect 52684 9976 52724 10016
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 55084 14428 55124 14468
rect 54700 14008 54740 14048
rect 55180 13252 55220 13292
rect 55372 13168 55412 13208
rect 55276 13084 55316 13124
rect 54604 13000 54644 13040
rect 54892 13000 54932 13040
rect 55564 15436 55604 15476
rect 55564 15268 55604 15308
rect 56044 14680 56084 14720
rect 56332 14680 56372 14720
rect 55948 14428 55988 14468
rect 56428 13840 56468 13880
rect 56524 13672 56564 13712
rect 56236 13588 56276 13628
rect 56140 13420 56180 13460
rect 56044 13168 56084 13208
rect 57945 17116 57985 17156
rect 57292 16444 57332 16484
rect 57292 16024 57332 16064
rect 57004 15268 57044 15308
rect 56908 14512 56948 14552
rect 56812 13504 56852 13544
rect 56332 13168 56372 13208
rect 56428 13084 56468 13124
rect 54412 12496 54452 12536
rect 55468 12496 55508 12536
rect 56140 12496 56180 12536
rect 56236 12160 56276 12200
rect 53356 11656 53396 11696
rect 53932 11656 53972 11696
rect 53356 10984 53396 11024
rect 53356 10732 53396 10772
rect 53740 11068 53780 11108
rect 52972 10144 53012 10184
rect 53836 10732 53876 10772
rect 53164 10060 53204 10100
rect 53644 10060 53684 10100
rect 53068 9892 53108 9932
rect 53068 9640 53108 9680
rect 52396 9556 52436 9596
rect 52204 8716 52244 8756
rect 52108 8632 52148 8672
rect 52396 8632 52436 8672
rect 53452 9976 53492 10016
rect 52684 9220 52724 9260
rect 52684 8884 52724 8924
rect 53260 8884 53300 8924
rect 52876 8800 52916 8840
rect 52780 8464 52820 8504
rect 53164 8632 53204 8672
rect 52972 8380 53012 8420
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 52204 8044 52244 8084
rect 52684 8044 52724 8084
rect 50092 6448 50132 6488
rect 50860 6448 50900 6488
rect 50380 6112 50420 6152
rect 49132 5608 49172 5648
rect 48940 5440 48980 5480
rect 49132 5104 49172 5144
rect 50380 5524 50420 5564
rect 49228 5020 49268 5060
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 49612 3592 49652 3632
rect 50668 4180 50708 4220
rect 50188 3592 50228 3632
rect 51724 6448 51764 6488
rect 51244 6196 51284 6236
rect 51436 6196 51476 6236
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 53932 10144 53972 10184
rect 53740 9472 53780 9512
rect 53452 8968 53492 9008
rect 53548 8884 53588 8924
rect 53452 8632 53492 8672
rect 53740 8800 53780 8840
rect 53356 8464 53396 8504
rect 53644 8380 53684 8420
rect 53260 8044 53300 8084
rect 52972 7792 53012 7832
rect 52876 7204 52916 7244
rect 53068 7120 53108 7160
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 52396 6196 52436 6236
rect 52012 5104 52052 5144
rect 52300 5608 52340 5648
rect 52780 5776 52820 5816
rect 52684 5692 52724 5732
rect 56236 11656 56276 11696
rect 56716 13168 56756 13208
rect 56908 13252 56948 13292
rect 56620 13000 56660 13040
rect 56812 11740 56852 11780
rect 54124 10984 54164 11024
rect 54028 8800 54068 8840
rect 54220 8968 54260 9008
rect 53932 8632 53972 8672
rect 53836 7960 53876 8000
rect 53452 7204 53492 7244
rect 53740 7204 53780 7244
rect 53356 7036 53396 7076
rect 53164 5776 53204 5816
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 52300 5104 52340 5144
rect 51820 5020 51860 5060
rect 51628 4768 51668 4808
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 51532 4348 51572 4388
rect 50860 4012 50900 4052
rect 50764 3928 50804 3968
rect 50860 3592 50900 3632
rect 51628 3424 51668 3464
rect 52108 4936 52148 4976
rect 52588 5020 52628 5060
rect 52492 4936 52532 4976
rect 52972 5608 53012 5648
rect 52300 4348 52340 4388
rect 51916 4264 51956 4304
rect 52684 4264 52724 4304
rect 53260 5020 53300 5060
rect 53068 4180 53108 4220
rect 52972 3928 53012 3968
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 52012 3592 52052 3632
rect 50092 3256 50132 3296
rect 51724 3256 51764 3296
rect 52684 3424 52724 3464
rect 52588 3256 52628 3296
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 3340 2584 3380 2624
rect 6028 2584 6068 2624
rect 54220 7960 54260 8000
rect 54508 9472 54548 9512
rect 54412 8800 54452 8840
rect 56428 10396 56468 10436
rect 55084 8548 55124 8588
rect 55660 8548 55700 8588
rect 55948 8548 55988 8588
rect 55180 8380 55220 8420
rect 54220 6532 54260 6572
rect 53548 5692 53588 5732
rect 53452 4936 53492 4976
rect 53548 4348 53588 4388
rect 53932 5608 53972 5648
rect 54220 5608 54260 5648
rect 54412 6448 54452 6488
rect 54700 7204 54740 7244
rect 54604 6532 54644 6572
rect 54796 6448 54836 6488
rect 54316 5524 54356 5564
rect 54124 5440 54164 5480
rect 54028 4768 54068 4808
rect 53836 3844 53876 3884
rect 53836 3508 53876 3548
rect 54700 5608 54740 5648
rect 54892 5524 54932 5564
rect 54892 4348 54932 4388
rect 54700 4264 54740 4304
rect 54604 4012 54644 4052
rect 54508 3424 54548 3464
rect 53740 2752 53780 2792
rect 53164 2500 53204 2540
rect 1036 2248 1076 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56812 8968 56852 9008
rect 57196 14848 57236 14888
rect 57100 13672 57140 13712
rect 58345 17200 58385 17240
rect 58540 16192 58580 16232
rect 58924 15772 58964 15812
rect 57484 14848 57524 14888
rect 57580 14680 57620 14720
rect 57676 14596 57716 14636
rect 57388 13420 57428 13460
rect 58348 14428 58388 14468
rect 57964 14260 58004 14300
rect 57772 14008 57812 14048
rect 58828 14512 58868 14552
rect 57868 13756 57908 13796
rect 57964 13504 58004 13544
rect 57676 13000 57716 13040
rect 57868 13000 57908 13040
rect 57292 12664 57332 12704
rect 57580 12496 57620 12536
rect 57484 11992 57524 12032
rect 57292 11572 57332 11612
rect 58348 13840 58388 13880
rect 58252 12664 58292 12704
rect 58060 12244 58100 12284
rect 58540 13168 58580 13208
rect 59020 13756 59060 13796
rect 58924 13168 58964 13208
rect 59500 15940 59540 15980
rect 59500 14680 59540 14720
rect 59500 14512 59540 14552
rect 59404 14344 59444 14384
rect 59308 12748 59348 12788
rect 59308 12580 59348 12620
rect 59020 12496 59060 12536
rect 58252 12244 58292 12284
rect 59116 12244 59156 12284
rect 59020 12076 59060 12116
rect 57964 11740 58004 11780
rect 58156 11740 58196 11780
rect 58348 11740 58388 11780
rect 58348 11572 58388 11612
rect 57580 10312 57620 10352
rect 57388 10228 57428 10268
rect 58060 10396 58100 10436
rect 57868 10144 57908 10184
rect 58444 11152 58484 11192
rect 58252 10312 58292 10352
rect 58060 9976 58100 10016
rect 57196 9136 57236 9176
rect 58348 9976 58388 10016
rect 58060 9052 58100 9092
rect 57772 8800 57812 8840
rect 57964 8800 58004 8840
rect 57868 8464 57908 8504
rect 56812 6280 56852 6320
rect 55852 5692 55892 5732
rect 56236 5524 56276 5564
rect 55660 4768 55700 4808
rect 55948 4936 55988 4976
rect 56332 4936 56372 4976
rect 56332 4768 56372 4808
rect 55852 4348 55892 4388
rect 55180 4264 55220 4304
rect 55660 4180 55700 4220
rect 55564 4096 55604 4136
rect 55084 3760 55124 3800
rect 55756 3928 55796 3968
rect 55948 3928 55988 3968
rect 55756 3760 55796 3800
rect 55468 2164 55508 2204
rect 53452 1744 53492 1784
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 56140 3844 56180 3884
rect 56140 3508 56180 3548
rect 55756 2752 55796 2792
rect 55852 2668 55892 2708
rect 56044 2500 56084 2540
rect 55852 2080 55892 2120
rect 56044 2164 56084 2204
rect 55948 1912 55988 1952
rect 55948 1744 55988 1784
rect 55756 1156 55796 1196
rect 56236 2752 56276 2792
rect 57772 6784 57812 6824
rect 57388 5692 57428 5732
rect 57004 5608 57044 5648
rect 56428 4684 56468 4724
rect 56716 4348 56756 4388
rect 57196 4348 57236 4388
rect 58348 9136 58388 9176
rect 58252 9052 58292 9092
rect 58252 8716 58292 8756
rect 58828 11656 58868 11696
rect 58924 11572 58964 11612
rect 58828 11152 58868 11192
rect 59404 12244 59444 12284
rect 59308 11572 59348 11612
rect 59308 11152 59348 11192
rect 59500 11488 59540 11528
rect 59692 12496 59732 12536
rect 58732 10228 58772 10268
rect 58636 9304 58676 9344
rect 58732 9052 58772 9092
rect 58540 8800 58580 8840
rect 58924 10228 58964 10268
rect 59212 10144 59252 10184
rect 59692 10984 59732 11024
rect 61545 17200 61585 17240
rect 61804 17200 61844 17240
rect 60172 16192 60212 16232
rect 60076 10816 60116 10856
rect 59884 10060 59924 10100
rect 59308 9220 59348 9260
rect 59212 9136 59252 9176
rect 59308 9052 59348 9092
rect 59020 8884 59060 8924
rect 59692 8884 59732 8924
rect 58444 8464 58484 8504
rect 58156 7960 58196 8000
rect 58732 8464 58772 8504
rect 57868 6364 57908 6404
rect 58060 6448 58100 6488
rect 58060 6280 58100 6320
rect 57964 5692 58004 5732
rect 58828 7960 58868 8000
rect 59404 8632 59444 8672
rect 59692 8716 59732 8756
rect 59308 8548 59348 8588
rect 59980 9976 60020 10016
rect 61708 16444 61748 16484
rect 61708 16276 61748 16316
rect 61612 16108 61652 16148
rect 61132 16024 61172 16064
rect 61420 16024 61460 16064
rect 62345 17200 62385 17240
rect 62188 16444 62228 16484
rect 61900 16192 61940 16232
rect 61804 15856 61844 15896
rect 62380 16192 62420 16232
rect 62668 17032 62708 17072
rect 62668 16108 62708 16148
rect 62092 15856 62132 15896
rect 61612 15268 61652 15308
rect 61612 14764 61652 14804
rect 60748 14680 60788 14720
rect 60460 14344 60500 14384
rect 60652 14260 60692 14300
rect 60556 13924 60596 13964
rect 61228 14680 61268 14720
rect 61996 15520 62036 15560
rect 62380 15268 62420 15308
rect 62284 14680 62324 14720
rect 61804 14512 61844 14552
rect 62188 14512 62228 14552
rect 61708 14344 61748 14384
rect 60844 14008 60884 14048
rect 60748 11824 60788 11864
rect 60748 11656 60788 11696
rect 62572 14428 62612 14468
rect 62476 14344 62516 14384
rect 61420 14092 61460 14132
rect 62380 14092 62420 14132
rect 61132 13000 61172 13040
rect 61324 13168 61364 13208
rect 62476 14008 62516 14048
rect 61708 13924 61748 13964
rect 61612 13336 61652 13376
rect 62572 13924 62612 13964
rect 62476 13336 62516 13376
rect 61996 13252 62036 13292
rect 61996 13000 62036 13040
rect 62284 13168 62324 13208
rect 61708 12580 61748 12620
rect 61612 12328 61652 12368
rect 61036 11908 61076 11948
rect 60844 11488 60884 11528
rect 60940 11152 60980 11192
rect 60364 10480 60404 10520
rect 60268 9976 60308 10016
rect 60844 9472 60884 9512
rect 59884 9052 59924 9092
rect 59308 8296 59348 8336
rect 59020 7960 59060 8000
rect 58924 7120 58964 7160
rect 58348 6616 58388 6656
rect 58828 6616 58868 6656
rect 58540 6448 58580 6488
rect 58252 6280 58292 6320
rect 58156 5524 58196 5564
rect 56524 3928 56564 3968
rect 56620 3424 56660 3464
rect 57004 4096 57044 4136
rect 57292 4264 57332 4304
rect 57964 4264 58004 4304
rect 58540 4684 58580 4724
rect 58828 6448 58868 6488
rect 58732 6364 58772 6404
rect 58828 5440 58868 5480
rect 59212 7036 59252 7076
rect 59020 6784 59060 6824
rect 59020 6616 59060 6656
rect 59692 7204 59732 7244
rect 59692 6700 59732 6740
rect 59212 6448 59252 6488
rect 59500 6448 59540 6488
rect 59020 6364 59060 6404
rect 58636 4180 58676 4220
rect 58252 4096 58292 4136
rect 58924 4096 58964 4136
rect 59404 5608 59444 5648
rect 59308 5440 59348 5480
rect 59212 4936 59252 4976
rect 59116 4180 59156 4220
rect 57100 3508 57140 3548
rect 58828 3424 58868 3464
rect 56524 2752 56564 2792
rect 59692 6532 59732 6572
rect 59788 6448 59828 6488
rect 59692 4936 59732 4976
rect 59404 4264 59444 4304
rect 59596 4264 59636 4304
rect 59500 3676 59540 3716
rect 59020 3088 59060 3128
rect 58924 2836 58964 2876
rect 56908 2752 56948 2792
rect 57292 2668 57332 2708
rect 58732 2668 58772 2708
rect 56524 2080 56564 2120
rect 56332 1912 56372 1952
rect 56524 1156 56564 1196
rect 57196 2080 57236 2120
rect 57004 1912 57044 1952
rect 57196 1408 57236 1448
rect 56428 1072 56468 1112
rect 57196 1072 57236 1112
rect 57580 2500 57620 2540
rect 57388 1912 57428 1952
rect 57868 1912 57908 1952
rect 57484 1072 57524 1112
rect 58636 1072 58676 1112
rect 59020 2668 59060 2708
rect 59404 3004 59444 3044
rect 59692 3424 59732 3464
rect 59788 2500 59828 2540
rect 59116 1912 59156 1952
rect 59020 1660 59060 1700
rect 59020 1408 59060 1448
rect 58924 1324 58964 1364
rect 59212 1324 59252 1364
rect 59596 1240 59636 1280
rect 60172 9220 60212 9260
rect 60076 8632 60116 8672
rect 60364 9136 60404 9176
rect 60268 8464 60308 8504
rect 59980 8296 60020 8336
rect 60076 8128 60116 8168
rect 60364 7792 60404 7832
rect 60172 7708 60212 7748
rect 60556 7708 60596 7748
rect 60460 7204 60500 7244
rect 60076 7036 60116 7076
rect 60172 6448 60212 6488
rect 60076 5692 60116 5732
rect 60268 6280 60308 6320
rect 62188 12916 62228 12956
rect 62092 12664 62132 12704
rect 61804 11404 61844 11444
rect 61804 10984 61844 11024
rect 62284 12412 62324 12452
rect 62092 12328 62132 12368
rect 62092 11656 62132 11696
rect 62572 11908 62612 11948
rect 62572 11740 62612 11780
rect 62380 11152 62420 11192
rect 62188 10984 62228 11024
rect 61996 10312 62036 10352
rect 61996 9640 62036 9680
rect 62188 9556 62228 9596
rect 61996 9220 62036 9260
rect 63532 16024 63572 16064
rect 64588 17116 64628 17156
rect 64855 17116 64895 17156
rect 62764 14848 62804 14888
rect 62956 15268 62996 15308
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 64684 16864 64724 16904
rect 65356 16528 65396 16568
rect 64972 16192 65012 16232
rect 64492 15688 64532 15728
rect 64780 15688 64820 15728
rect 64108 15352 64148 15392
rect 63820 14680 63860 14720
rect 64972 15520 65012 15560
rect 64684 14680 64724 14720
rect 66604 17116 66644 17156
rect 66855 17116 66895 17156
rect 66796 16192 66836 16232
rect 66124 15940 66164 15980
rect 65740 15268 65780 15308
rect 66220 15436 66260 15476
rect 63916 14512 63956 14552
rect 63724 14344 63764 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 63916 13924 63956 13964
rect 63532 13420 63572 13460
rect 62860 13252 62900 13292
rect 64396 13924 64436 13964
rect 64108 13336 64148 13376
rect 63628 13168 63668 13208
rect 63916 13168 63956 13208
rect 62860 13084 62900 13124
rect 62764 12160 62804 12200
rect 62764 11908 62804 11948
rect 63820 13000 63860 13040
rect 63532 12916 63572 12956
rect 64012 12916 64052 12956
rect 63340 12496 63380 12536
rect 63244 12328 63284 12368
rect 63052 12244 63092 12284
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 64396 13336 64436 13376
rect 64588 13000 64628 13040
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 64204 12664 64244 12704
rect 64396 12496 64436 12536
rect 63724 12412 63764 12452
rect 63628 12244 63668 12284
rect 62764 11572 62804 11612
rect 63244 11908 63284 11948
rect 63532 11908 63572 11948
rect 63436 11824 63476 11864
rect 63436 11404 63476 11444
rect 63244 11320 63284 11360
rect 62764 11152 62804 11192
rect 62668 8968 62708 9008
rect 64588 12412 64628 12452
rect 64012 12328 64052 12368
rect 63820 11572 63860 11612
rect 63916 11404 63956 11444
rect 63820 11320 63860 11360
rect 62956 10984 62996 11024
rect 63916 10984 63956 11024
rect 64204 11824 64244 11864
rect 64396 12076 64436 12116
rect 65164 14680 65204 14720
rect 65932 14008 65972 14048
rect 65548 13840 65588 13880
rect 64876 11824 64916 11864
rect 65548 12496 65588 12536
rect 66028 12496 66068 12536
rect 64588 11740 64628 11780
rect 64972 11740 65012 11780
rect 65452 11740 65492 11780
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 63436 10396 63476 10436
rect 63436 10144 63476 10184
rect 63628 10060 63668 10100
rect 63436 9472 63476 9512
rect 63820 9220 63860 9260
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 62860 8800 62900 8840
rect 62860 8632 62900 8672
rect 64204 10144 64244 10184
rect 64588 10984 64628 11024
rect 64684 10900 64724 10940
rect 64588 10396 64628 10436
rect 65164 10900 65204 10940
rect 64108 8968 64148 9008
rect 64012 8632 64052 8672
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 64876 9556 64916 9596
rect 64588 9220 64628 9260
rect 65164 10060 65204 10100
rect 64780 8968 64820 9008
rect 64396 8800 64436 8840
rect 65068 8800 65108 8840
rect 65452 10396 65492 10436
rect 66508 14260 66548 14300
rect 66700 14008 66740 14048
rect 66220 11992 66260 12032
rect 66028 11656 66068 11696
rect 67372 16192 67412 16232
rect 67276 16108 67316 16148
rect 67180 14764 67220 14804
rect 67564 14596 67604 14636
rect 66988 14260 67028 14300
rect 66892 12580 66932 12620
rect 66892 10060 66932 10100
rect 66796 9640 66836 9680
rect 66604 9472 66644 9512
rect 64492 8464 64532 8504
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 62860 8128 62900 8168
rect 60844 7120 60884 7160
rect 60652 6280 60692 6320
rect 61036 7120 61076 7160
rect 64876 8464 64916 8504
rect 63820 7960 63860 8000
rect 62188 7708 62228 7748
rect 63628 7708 63668 7748
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 61324 6448 61364 6488
rect 61900 6448 61940 6488
rect 60940 6112 60980 6152
rect 60652 5692 60692 5732
rect 60172 5020 60212 5060
rect 60076 4936 60116 4976
rect 59980 4180 60020 4220
rect 60460 5020 60500 5060
rect 60364 3004 60404 3044
rect 59980 2920 60020 2960
rect 60364 2668 60404 2708
rect 61324 5608 61364 5648
rect 61516 5608 61556 5648
rect 61036 5104 61076 5144
rect 60940 4936 60980 4976
rect 60748 4096 60788 4136
rect 61420 5104 61460 5144
rect 61612 5020 61652 5060
rect 63436 6196 63476 6236
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 63340 5860 63380 5900
rect 61996 5692 62036 5732
rect 61516 4936 61556 4976
rect 61612 4852 61652 4892
rect 62476 5608 62516 5648
rect 62956 5440 62996 5480
rect 64108 7120 64148 7160
rect 63916 7036 63956 7076
rect 63916 6700 63956 6740
rect 63628 5692 63668 5732
rect 63532 5608 63572 5648
rect 63628 5524 63668 5564
rect 64108 6448 64148 6488
rect 64396 7960 64436 8000
rect 64780 7960 64820 8000
rect 64684 7792 64724 7832
rect 65068 7960 65108 8000
rect 65548 7960 65588 8000
rect 65260 7876 65300 7916
rect 65164 7708 65204 7748
rect 65740 7876 65780 7916
rect 65644 7792 65684 7832
rect 64300 7120 64340 7160
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 64972 7120 65012 7160
rect 64876 7036 64916 7076
rect 64780 6700 64820 6740
rect 65260 6868 65300 6908
rect 65548 6868 65588 6908
rect 65260 6448 65300 6488
rect 64204 5776 64244 5816
rect 63628 4936 63668 4976
rect 63916 4936 63956 4976
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 61804 4264 61844 4304
rect 62764 4264 62804 4304
rect 61228 4096 61268 4136
rect 60556 3088 60596 3128
rect 60460 1912 60500 1952
rect 59884 1072 59924 1112
rect 60076 1072 60116 1112
rect 60652 2500 60692 2540
rect 60556 1156 60596 1196
rect 62092 3676 62132 3716
rect 62860 3592 62900 3632
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 62764 2920 62804 2960
rect 61612 2500 61652 2540
rect 60940 1912 60980 1952
rect 60844 1240 60884 1280
rect 61804 1324 61844 1364
rect 62476 1324 62516 1364
rect 62284 1240 62324 1280
rect 64588 5776 64628 5816
rect 65068 5776 65108 5816
rect 64204 5608 64244 5648
rect 64780 5608 64820 5648
rect 64684 5440 64724 5480
rect 64780 5356 64820 5396
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 64012 4264 64052 4304
rect 64012 3592 64052 3632
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 65164 5692 65204 5732
rect 65356 6280 65396 6320
rect 65260 5356 65300 5396
rect 64876 5104 64916 5144
rect 66604 8632 66644 8672
rect 67084 13924 67124 13964
rect 67276 13924 67316 13964
rect 67372 13840 67412 13880
rect 67564 13840 67604 13880
rect 67468 13252 67508 13292
rect 67948 16192 67988 16232
rect 67852 15688 67892 15728
rect 68524 16024 68564 16064
rect 69004 16192 69044 16232
rect 69388 16108 69428 16148
rect 70156 16192 70196 16232
rect 71404 17116 71444 17156
rect 71655 17116 71695 17156
rect 70527 16024 70567 16064
rect 69100 15940 69140 15980
rect 69772 15940 69812 15980
rect 68716 15436 68756 15476
rect 68236 14596 68276 14636
rect 67852 13672 67892 13712
rect 67180 12748 67220 12788
rect 67180 12412 67220 12452
rect 67372 11572 67412 11612
rect 67276 10312 67316 10352
rect 67276 8632 67316 8672
rect 66028 7708 66068 7748
rect 65740 7120 65780 7160
rect 65836 7121 65876 7160
rect 65836 7120 65876 7121
rect 65548 5440 65588 5480
rect 65164 5020 65204 5060
rect 63916 3424 63956 3464
rect 64588 3424 64628 3464
rect 64108 3256 64148 3296
rect 63052 1912 63092 1952
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 62860 1156 62900 1196
rect 61996 988 62036 1028
rect 63628 988 63668 1028
rect 63820 2416 63860 2456
rect 65644 5104 65684 5144
rect 66220 6868 66260 6908
rect 65932 6448 65972 6488
rect 65836 6280 65876 6320
rect 66604 7120 66644 7160
rect 66220 5608 66260 5648
rect 66508 5608 66548 5648
rect 66796 7036 66836 7076
rect 66796 6448 66836 6488
rect 66124 5440 66164 5480
rect 66316 5440 66356 5480
rect 66124 5020 66164 5060
rect 65548 4936 65588 4976
rect 65740 4936 65780 4976
rect 65260 4012 65300 4052
rect 65260 3424 65300 3464
rect 65452 3256 65492 3296
rect 64204 2836 64244 2876
rect 64492 2668 64532 2708
rect 64780 2668 64820 2708
rect 64396 2500 64436 2540
rect 64780 2500 64820 2540
rect 64684 2416 64724 2456
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 64108 1408 64148 1448
rect 65164 2080 65204 2120
rect 64780 1240 64820 1280
rect 65164 1408 65204 1448
rect 65836 4264 65876 4304
rect 65932 4012 65972 4052
rect 66508 4936 66548 4976
rect 66028 3340 66068 3380
rect 66700 4432 66740 4472
rect 66316 3340 66356 3380
rect 67660 10396 67700 10436
rect 67852 10312 67892 10352
rect 67756 8128 67796 8168
rect 67852 7120 67892 7160
rect 68332 14344 68372 14384
rect 68524 14344 68564 14384
rect 68140 13924 68180 13964
rect 68044 13840 68084 13880
rect 68140 13756 68180 13796
rect 68044 13672 68084 13712
rect 67948 5524 67988 5564
rect 67756 4684 67796 4724
rect 67372 3676 67412 3716
rect 66124 2836 66164 2876
rect 65740 2416 65780 2456
rect 65740 1912 65780 1952
rect 66028 1156 66068 1196
rect 67372 2416 67412 2456
rect 66892 2080 66932 2120
rect 67276 1912 67316 1952
rect 67468 1912 67508 1952
rect 67948 2248 67988 2288
rect 67564 1828 67604 1868
rect 68812 14092 68852 14132
rect 69868 15352 69908 15392
rect 69196 14344 69236 14384
rect 69100 14260 69140 14300
rect 69388 14092 69428 14132
rect 68524 13588 68564 13628
rect 68716 13588 68756 13628
rect 68428 13420 68468 13460
rect 68812 13420 68852 13460
rect 68620 13000 68660 13040
rect 68620 12832 68660 12872
rect 68620 12496 68660 12536
rect 68908 13168 68948 13208
rect 69196 13840 69236 13880
rect 69292 13756 69332 13796
rect 69100 13588 69140 13628
rect 69100 13252 69140 13292
rect 69004 12916 69044 12956
rect 69100 12496 69140 12536
rect 68812 11824 68852 11864
rect 69004 11824 69044 11864
rect 68908 11656 68948 11696
rect 69868 15016 69908 15056
rect 70156 14428 70196 14468
rect 70060 14092 70100 14132
rect 69964 14008 70004 14048
rect 69868 13924 69908 13964
rect 70732 15520 70772 15560
rect 70540 15268 70580 15308
rect 70636 14932 70676 14972
rect 70828 15100 70868 15140
rect 70732 14848 70772 14888
rect 70636 14680 70676 14720
rect 70540 14512 70580 14552
rect 69868 13504 69908 13544
rect 70156 13504 70196 13544
rect 69580 13168 69620 13208
rect 69484 13000 69524 13040
rect 69484 11908 69524 11948
rect 69292 11656 69332 11696
rect 69004 11572 69044 11612
rect 69772 12832 69812 12872
rect 69676 12076 69716 12116
rect 70156 13000 70196 13040
rect 70060 12832 70100 12872
rect 70060 12496 70100 12536
rect 69964 11992 70004 12032
rect 69868 11908 69908 11948
rect 70060 11824 70100 11864
rect 69868 11740 69908 11780
rect 69676 11068 69716 11108
rect 68908 10564 68948 10604
rect 68428 10480 68468 10520
rect 68236 10228 68276 10268
rect 68908 10312 68948 10352
rect 68620 10228 68660 10268
rect 68524 10144 68564 10184
rect 70828 14512 70868 14552
rect 71116 15268 71156 15308
rect 71308 15100 71348 15140
rect 71020 14428 71060 14468
rect 71116 14008 71156 14048
rect 70924 13840 70964 13880
rect 70828 13756 70868 13796
rect 70636 12664 70676 12704
rect 70252 12496 70292 12536
rect 70252 12160 70292 12200
rect 70348 12076 70388 12116
rect 70252 11572 70292 11612
rect 70156 11068 70196 11108
rect 70540 11992 70580 12032
rect 70636 11740 70676 11780
rect 70444 11656 70484 11696
rect 70348 11236 70388 11276
rect 69388 10564 69428 10604
rect 69292 10228 69332 10268
rect 69196 10144 69236 10184
rect 68812 10060 68852 10100
rect 69100 10060 69140 10100
rect 68332 9892 68372 9932
rect 68140 8632 68180 8672
rect 68140 7120 68180 7160
rect 68908 9220 68948 9260
rect 68428 8296 68468 8336
rect 68716 8632 68756 8672
rect 69004 8800 69044 8840
rect 68428 7708 68468 7748
rect 69484 10480 69524 10520
rect 69772 10312 69812 10352
rect 69676 10144 69716 10184
rect 69580 10060 69620 10100
rect 69676 9892 69716 9932
rect 69388 9388 69428 9428
rect 69292 8968 69332 9008
rect 69196 8800 69236 8840
rect 69196 8548 69236 8588
rect 69388 8800 69428 8840
rect 69676 8968 69716 9008
rect 69868 9556 69908 9596
rect 69868 9304 69908 9344
rect 69580 8632 69620 8672
rect 69100 7036 69140 7076
rect 69676 8464 69716 8504
rect 69388 6028 69428 6068
rect 69196 5860 69236 5900
rect 69100 5608 69140 5648
rect 69292 5627 69332 5648
rect 69292 5608 69332 5627
rect 68236 4768 68276 4808
rect 68812 4684 68852 4724
rect 68812 4432 68852 4472
rect 68716 4264 68756 4304
rect 68236 3256 68276 3296
rect 68812 4096 68852 4136
rect 68716 3088 68756 3128
rect 68332 2500 68372 2540
rect 68140 2416 68180 2456
rect 68236 2332 68276 2372
rect 68044 1660 68084 1700
rect 68524 1828 68564 1868
rect 67372 1156 67412 1196
rect 58924 904 58964 944
rect 60364 904 60404 944
rect 62956 904 62996 944
rect 63724 904 63764 944
rect 64204 904 64244 944
rect 70060 10312 70100 10352
rect 70156 9472 70196 9512
rect 70156 8800 70196 8840
rect 70060 8548 70100 8588
rect 69868 7204 69908 7244
rect 69964 7120 70004 7160
rect 70732 10732 70772 10772
rect 71116 10732 71156 10772
rect 70636 10228 70676 10268
rect 70444 9304 70484 9344
rect 70540 9052 70580 9092
rect 70828 10144 70868 10184
rect 70924 9976 70964 10016
rect 70828 9472 70868 9512
rect 71308 10144 71348 10184
rect 71116 9892 71156 9932
rect 71596 12916 71636 12956
rect 71980 16108 72020 16148
rect 72556 15688 72596 15728
rect 72172 15184 72212 15224
rect 72172 14512 72212 14552
rect 72748 14008 72788 14048
rect 71788 12748 71828 12788
rect 71500 10396 71540 10436
rect 71692 10144 71732 10184
rect 71692 9892 71732 9932
rect 70732 8800 70772 8840
rect 70348 8464 70388 8504
rect 70348 7708 70388 7748
rect 70156 7120 70196 7160
rect 70348 7204 70388 7244
rect 69964 6448 70004 6488
rect 69772 6028 69812 6068
rect 69772 5860 69812 5900
rect 69196 4684 69236 4724
rect 69004 4264 69044 4304
rect 69004 3592 69044 3632
rect 68908 3424 68948 3464
rect 69292 3592 69332 3632
rect 69964 5608 70004 5648
rect 70540 7120 70580 7160
rect 70444 6448 70484 6488
rect 70444 4348 70484 4388
rect 70252 4264 70292 4304
rect 69964 3508 70004 3548
rect 69772 3256 69812 3296
rect 69004 3088 69044 3128
rect 70444 4096 70484 4136
rect 70252 3424 70292 3464
rect 69868 2500 69908 2540
rect 69196 2332 69236 2372
rect 71212 9556 71252 9596
rect 71116 9472 71156 9512
rect 71404 9220 71444 9260
rect 71308 9136 71348 9176
rect 71884 9472 71924 9512
rect 71692 9388 71732 9428
rect 71020 8296 71060 8336
rect 71020 7708 71060 7748
rect 71884 9220 71924 9260
rect 72172 13168 72212 13208
rect 73036 12916 73076 12956
rect 72844 12664 72884 12704
rect 72460 11152 72500 11192
rect 72844 10396 72884 10436
rect 72940 10144 72980 10184
rect 72844 10060 72884 10100
rect 72556 9724 72596 9764
rect 72556 9388 72596 9428
rect 70828 5608 70868 5648
rect 71308 5608 71348 5648
rect 71788 6784 71828 6824
rect 71980 7120 72020 7160
rect 71980 6784 72020 6824
rect 71692 5692 71732 5732
rect 71596 5608 71636 5648
rect 71884 6448 71924 6488
rect 71980 5776 72020 5816
rect 71788 5524 71828 5564
rect 70828 4936 70868 4976
rect 70636 4348 70676 4388
rect 70732 4264 70772 4304
rect 70732 3592 70772 3632
rect 70636 3508 70676 3548
rect 70540 3340 70580 3380
rect 69004 1828 69044 1868
rect 70060 1912 70100 1952
rect 70252 1912 70292 1952
rect 70924 3340 70964 3380
rect 71308 4684 71348 4724
rect 71500 4936 71540 4976
rect 71884 4936 71924 4976
rect 71788 4852 71828 4892
rect 71404 4348 71444 4388
rect 71308 4264 71348 4304
rect 71020 2668 71060 2708
rect 71212 2836 71252 2876
rect 71788 3676 71828 3716
rect 71404 3508 71444 3548
rect 71596 3508 71636 3548
rect 71692 3256 71732 3296
rect 71692 3088 71732 3128
rect 71884 2752 71924 2792
rect 71308 2668 71348 2708
rect 71788 2668 71828 2708
rect 71020 2332 71060 2372
rect 71212 2332 71252 2372
rect 70924 1912 70964 1952
rect 71788 1912 71828 1952
rect 70828 1828 70868 1868
rect 72172 5692 72212 5732
rect 72652 7120 72692 7160
rect 72940 6448 72980 6488
rect 72268 5524 72308 5564
rect 72172 4936 72212 4976
rect 72076 4264 72116 4304
rect 72076 3592 72116 3632
rect 72748 5608 72788 5648
rect 73420 12916 73460 12956
rect 73324 12664 73364 12704
rect 74284 15436 74324 15476
rect 73804 15268 73844 15308
rect 73612 14848 73652 14888
rect 74092 14848 74132 14888
rect 73708 14512 73748 14552
rect 73612 14428 73652 14468
rect 73516 10396 73556 10436
rect 73420 10060 73460 10100
rect 73516 7960 73556 8000
rect 74380 14596 74420 14636
rect 74188 14344 74228 14384
rect 74380 14344 74420 14384
rect 73900 13672 73940 13712
rect 73708 12916 73748 12956
rect 73996 12580 74036 12620
rect 73996 11740 74036 11780
rect 74860 16192 74900 16232
rect 75945 17200 75985 17240
rect 74668 15352 74708 15392
rect 74764 14764 74804 14804
rect 74668 14008 74708 14048
rect 75340 16192 75380 16232
rect 75724 16192 75764 16232
rect 74956 16108 74996 16148
rect 76588 16024 76628 16064
rect 77164 16192 77204 16232
rect 76972 15772 77012 15812
rect 75148 15520 75188 15560
rect 75244 15268 75284 15308
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 75628 15268 75668 15308
rect 75628 14848 75668 14888
rect 75628 14680 75668 14720
rect 75052 14596 75092 14636
rect 74956 14512 74996 14552
rect 75820 14680 75860 14720
rect 74860 14428 74900 14468
rect 76012 14512 76052 14552
rect 78988 17116 79028 17156
rect 74092 9472 74132 9512
rect 74956 13924 74996 13964
rect 74860 13840 74900 13880
rect 74764 13672 74804 13712
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 77164 14176 77204 14216
rect 75820 13756 75860 13796
rect 74860 13504 74900 13544
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 75148 13420 75188 13460
rect 74380 13336 74420 13376
rect 74572 13336 74612 13376
rect 74956 13336 74996 13376
rect 74284 13168 74324 13208
rect 74764 13168 74804 13208
rect 75052 13168 75092 13208
rect 74956 13084 74996 13124
rect 75724 13252 75764 13292
rect 75148 13084 75188 13124
rect 75820 13168 75860 13208
rect 75532 13000 75572 13040
rect 74476 12664 74516 12704
rect 74572 12328 74612 12368
rect 74764 12580 74804 12620
rect 74764 12328 74804 12368
rect 74668 10984 74708 11024
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 74956 11908 74996 11948
rect 74860 11320 74900 11360
rect 74668 10144 74708 10184
rect 74572 9556 74612 9596
rect 76492 13168 76532 13208
rect 77164 13252 77204 13292
rect 76972 13084 77012 13124
rect 76108 12664 76148 12704
rect 75820 12580 75860 12620
rect 75724 11908 75764 11948
rect 75628 11656 75668 11696
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 76780 12664 76820 12704
rect 76396 12496 76436 12536
rect 76876 12496 76916 12536
rect 75436 11488 75476 11528
rect 76012 11488 76052 11528
rect 75340 11320 75380 11360
rect 75244 11152 75284 11192
rect 75148 10984 75188 11024
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 75820 10984 75860 11024
rect 75916 10396 75956 10436
rect 74860 9640 74900 9680
rect 76204 11656 76244 11696
rect 77644 14008 77684 14048
rect 78220 14008 78260 14048
rect 76588 11656 76628 11696
rect 77068 11740 77108 11780
rect 76396 11572 76436 11612
rect 76300 11488 76340 11528
rect 77164 11572 77204 11612
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 76300 11152 76340 11192
rect 75916 10060 75956 10100
rect 75532 9808 75572 9848
rect 75724 9640 75764 9680
rect 75628 9556 75668 9596
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 76012 9808 76052 9848
rect 76684 10984 76724 11024
rect 76300 10060 76340 10100
rect 76588 10396 76628 10436
rect 76492 10228 76532 10268
rect 76396 9976 76436 10016
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 76492 9640 76532 9680
rect 75820 9220 75860 9260
rect 76204 9485 76244 9512
rect 76204 9472 76244 9485
rect 75724 8548 75764 8588
rect 74860 8044 74900 8084
rect 73228 6448 73268 6488
rect 73612 6448 73652 6488
rect 72460 4348 72500 4388
rect 72268 3508 72308 3548
rect 72460 3424 72500 3464
rect 72844 4348 72884 4388
rect 72748 3424 72788 3464
rect 75532 7960 75572 8000
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 75628 7876 75668 7916
rect 75436 7204 75476 7244
rect 75724 7792 75764 7832
rect 76588 9556 76628 9596
rect 77260 11152 77300 11192
rect 76876 10060 76916 10100
rect 76780 9388 76820 9428
rect 76684 9220 76724 9260
rect 77644 12916 77684 12956
rect 77644 12496 77684 12536
rect 78124 12496 78164 12536
rect 78412 15772 78452 15812
rect 78316 12244 78356 12284
rect 78316 11740 78356 11780
rect 77740 10228 77780 10268
rect 77356 9640 77396 9680
rect 76300 8548 76340 8588
rect 75916 8464 75956 8504
rect 75916 8128 75956 8168
rect 76588 8548 76628 8588
rect 76204 8380 76244 8420
rect 76108 7960 76148 8000
rect 75820 7288 75860 7328
rect 75724 7120 75764 7160
rect 75820 7036 75860 7076
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 76396 8128 76436 8168
rect 76300 8044 76340 8084
rect 76012 7792 76052 7832
rect 76204 7372 76244 7412
rect 77260 9472 77300 9512
rect 77548 9472 77588 9512
rect 78316 10144 78356 10184
rect 78124 9640 78164 9680
rect 77932 9472 77972 9512
rect 77356 9136 77396 9176
rect 76204 7204 76244 7244
rect 76588 7204 76628 7244
rect 74860 6532 74900 6572
rect 74764 6280 74804 6320
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 74380 5608 74420 5648
rect 74476 4768 74516 4808
rect 73708 4264 73748 4304
rect 74284 4264 74324 4304
rect 74476 4180 74516 4220
rect 75820 6784 75860 6824
rect 75724 6532 75764 6572
rect 75628 6448 75668 6488
rect 76108 7036 76148 7076
rect 76684 7120 76724 7160
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 76492 6532 76532 6572
rect 75628 6280 75668 6320
rect 76300 6448 76340 6488
rect 76588 6448 76628 6488
rect 76396 5608 76436 5648
rect 77260 7960 77300 8000
rect 78028 7960 78068 8000
rect 77164 7204 77204 7244
rect 77356 7288 77396 7328
rect 77260 7120 77300 7160
rect 77836 7288 77876 7328
rect 77644 7120 77684 7160
rect 77260 5608 77300 5648
rect 77644 6532 77684 6572
rect 76492 5440 76532 5480
rect 74860 4768 74900 4808
rect 74572 4096 74612 4136
rect 74764 4096 74804 4136
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 76108 5272 76148 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 76204 4348 76244 4388
rect 75820 4264 75860 4304
rect 75724 4096 75764 4136
rect 73708 3508 73748 3548
rect 76588 4936 76628 4976
rect 76396 4180 76436 4220
rect 76876 4264 76916 4304
rect 76780 4096 76820 4136
rect 76012 3592 76052 3632
rect 75820 3508 75860 3548
rect 72076 2668 72116 2708
rect 72172 2584 72212 2624
rect 72076 2416 72116 2456
rect 70732 1072 70772 1112
rect 71212 1072 71252 1112
rect 72844 3172 72884 3212
rect 73132 3424 73172 3464
rect 74572 3424 74612 3464
rect 73996 3256 74036 3296
rect 72940 2836 72980 2876
rect 73612 2752 73652 2792
rect 73900 2752 73940 2792
rect 72940 2668 72980 2708
rect 73708 2584 73748 2624
rect 73804 1912 73844 1952
rect 73228 1072 73268 1112
rect 74188 2668 74228 2708
rect 74476 2668 74516 2708
rect 73996 2500 74036 2540
rect 73996 2164 74036 2204
rect 74284 2584 74324 2624
rect 74476 2248 74516 2288
rect 74860 3340 74900 3380
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 74860 2920 74900 2960
rect 74668 2752 74708 2792
rect 74764 2584 74804 2624
rect 74668 2248 74708 2288
rect 73996 1828 74036 1868
rect 73996 1072 74036 1112
rect 74572 1912 74612 1952
rect 76108 3424 76148 3464
rect 76012 3088 76052 3128
rect 75820 2416 75860 2456
rect 75244 1912 75284 1952
rect 74764 1576 74804 1616
rect 75628 1576 75668 1616
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 76108 2920 76148 2960
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 76300 3592 76340 3632
rect 76780 3508 76820 3548
rect 76684 3424 76724 3464
rect 76396 3256 76436 3296
rect 76780 3256 76820 3296
rect 76396 2668 76436 2708
rect 76876 2920 76916 2960
rect 76108 2416 76148 2456
rect 76780 2416 76820 2456
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 77356 4936 77396 4976
rect 77452 4768 77492 4808
rect 77836 4768 77876 4808
rect 78604 14932 78644 14972
rect 78604 14512 78644 14552
rect 78892 16192 78932 16232
rect 79372 17116 79412 17156
rect 79655 17116 79695 17156
rect 79180 14932 79220 14972
rect 78700 14176 78740 14216
rect 79372 14176 79412 14216
rect 79276 12244 79316 12284
rect 79468 10228 79508 10268
rect 79468 9640 79508 9680
rect 79468 6532 79508 6572
rect 77836 4264 77876 4304
rect 78412 4264 78452 4304
rect 79468 4264 79508 4304
rect 77452 3172 77492 3212
rect 77836 3424 77876 3464
rect 77836 3172 77876 3212
rect 77356 2668 77396 2708
rect 77068 2584 77108 2624
rect 76972 2164 77012 2204
rect 78124 2920 78164 2960
rect 78316 2920 78356 2960
rect 77164 2416 77204 2456
rect 77356 2416 77396 2456
rect 77740 1912 77780 1952
rect 76204 1072 76244 1112
rect 76780 1072 76820 1112
rect 78028 1072 78068 1112
rect 78220 2164 78260 2204
rect 78220 1240 78260 1280
rect 78892 2584 78932 2624
rect 78700 2416 78740 2456
rect 78412 1912 78452 1952
rect 79468 1240 79508 1280
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 16343 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 16729 38576
rect 28343 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 28729 38576
rect 40343 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 40729 38576
rect 52343 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 52729 38576
rect 64343 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 64729 38576
rect 76343 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 76729 38576
rect 63340 38284 70156 38324
rect 70196 38284 71404 38324
rect 71444 38284 71453 38324
rect 59395 38240 59453 38241
rect 63340 38240 63380 38284
rect 59310 38200 59404 38240
rect 59444 38200 63380 38240
rect 67459 38200 67468 38240
rect 67508 38200 67517 38240
rect 59395 38199 59453 38200
rect 67468 38156 67508 38200
rect 57859 38116 57868 38156
rect 57908 38116 60020 38156
rect 67468 38116 69388 38156
rect 69428 38116 69437 38156
rect 59980 38072 60020 38116
rect 57283 38032 57292 38072
rect 57332 38032 59828 38072
rect 59971 38032 59980 38072
rect 60020 38032 60460 38072
rect 60500 38032 67756 38072
rect 67796 38032 67805 38072
rect 59788 37988 59828 38032
rect 55939 37948 55948 37988
rect 55988 37948 58060 37988
rect 58100 37948 58109 37988
rect 59779 37948 59788 37988
rect 59828 37948 61132 37988
rect 61172 37948 61181 37988
rect 63523 37948 63532 37988
rect 63572 37948 64300 37988
rect 64340 37948 64349 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 15103 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 15489 37820
rect 27103 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 27489 37820
rect 39103 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 39489 37820
rect 51103 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 51489 37820
rect 63103 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 63489 37820
rect 68707 37780 68716 37820
rect 68756 37780 69388 37820
rect 69428 37780 69437 37820
rect 75103 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 75489 37820
rect 67747 37612 67756 37652
rect 67796 37612 68236 37652
rect 68276 37612 68285 37652
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 0 37508 80 37528
rect 58339 37444 58348 37484
rect 58388 37444 60268 37484
rect 60308 37444 60317 37484
rect 73027 37444 73036 37484
rect 73076 37444 73612 37484
rect 73652 37444 73661 37484
rect 72451 37400 72509 37401
rect 76963 37400 77021 37401
rect 55363 37360 55372 37400
rect 55412 37360 55660 37400
rect 55700 37360 55709 37400
rect 57187 37360 57196 37400
rect 57236 37360 58828 37400
rect 58868 37360 58877 37400
rect 60355 37360 60364 37400
rect 60404 37360 62956 37400
rect 62996 37360 65548 37400
rect 65588 37360 65597 37400
rect 66307 37360 66316 37400
rect 66356 37360 67276 37400
rect 67316 37360 67325 37400
rect 72451 37360 72460 37400
rect 72500 37360 73228 37400
rect 73268 37360 73277 37400
rect 73987 37360 73996 37400
rect 74036 37360 74324 37400
rect 74755 37360 74764 37400
rect 74804 37360 76780 37400
rect 76820 37360 76829 37400
rect 76963 37360 76972 37400
rect 77012 37360 77164 37400
rect 77204 37360 77213 37400
rect 77443 37360 77452 37400
rect 77492 37360 78508 37400
rect 78548 37360 78557 37400
rect 57196 37232 57236 37360
rect 72451 37359 72509 37360
rect 74284 37316 74324 37360
rect 76963 37359 77021 37360
rect 77164 37316 77204 37360
rect 57475 37276 57484 37316
rect 57524 37276 58060 37316
rect 58100 37276 58732 37316
rect 58772 37276 61612 37316
rect 61652 37276 61661 37316
rect 63427 37276 63436 37316
rect 63476 37276 64204 37316
rect 64244 37276 66700 37316
rect 66740 37276 66749 37316
rect 67939 37276 67948 37316
rect 67988 37276 68140 37316
rect 68180 37276 68428 37316
rect 68468 37276 68477 37316
rect 73411 37276 73420 37316
rect 73460 37276 73900 37316
rect 73940 37276 74132 37316
rect 74284 37276 74380 37316
rect 74420 37276 74429 37316
rect 77164 37276 78316 37316
rect 78356 37276 79468 37316
rect 79508 37276 79517 37316
rect 55651 37192 55660 37232
rect 55700 37192 56716 37232
rect 56756 37192 57236 37232
rect 58147 37192 58156 37232
rect 58196 37192 58828 37232
rect 58868 37192 58877 37232
rect 63523 37192 63532 37232
rect 63572 37192 64108 37232
rect 64148 37192 64157 37232
rect 68323 37192 68332 37232
rect 68372 37192 69484 37232
rect 69524 37192 69533 37232
rect 71107 37192 71116 37232
rect 71156 37192 71500 37232
rect 71540 37192 71549 37232
rect 72931 37192 72940 37232
rect 72980 37192 72989 37232
rect 72940 37148 72980 37192
rect 67555 37108 67564 37148
rect 67604 37108 74036 37148
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 16343 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 16729 37064
rect 28343 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 28729 37064
rect 40343 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 40729 37064
rect 52343 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 52729 37064
rect 64343 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 64729 37064
rect 71971 37024 71980 37064
rect 72020 37024 72940 37064
rect 72980 37024 72989 37064
rect 58531 36940 58540 36980
rect 58580 36940 59788 36980
rect 59828 36940 61516 36980
rect 61556 36940 69196 36980
rect 69236 36940 69245 36980
rect 69091 36896 69149 36897
rect 73996 36896 74036 37108
rect 74092 36980 74132 37276
rect 74563 37192 74572 37232
rect 74612 37192 75052 37232
rect 75092 37192 77260 37232
rect 77300 37192 77932 37232
rect 77972 37192 77981 37232
rect 76343 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 76729 37064
rect 74083 36940 74092 36980
rect 74132 36940 74141 36980
rect 55747 36856 55756 36896
rect 55796 36856 57100 36896
rect 57140 36856 57149 36896
rect 58243 36856 58252 36896
rect 58292 36856 59020 36896
rect 59060 36856 59308 36896
rect 59348 36856 59357 36896
rect 67363 36856 67372 36896
rect 67412 36856 68140 36896
rect 68180 36856 68189 36896
rect 69006 36856 69100 36896
rect 69140 36856 69149 36896
rect 69283 36856 69292 36896
rect 69332 36856 70540 36896
rect 70580 36856 70589 36896
rect 73219 36856 73228 36896
rect 73268 36856 73940 36896
rect 73996 36856 75244 36896
rect 75284 36856 75293 36896
rect 69091 36855 69149 36856
rect 73900 36812 73940 36856
rect 54403 36772 54412 36812
rect 54452 36772 55564 36812
rect 55604 36772 55613 36812
rect 69475 36772 69484 36812
rect 69524 36772 71116 36812
rect 71156 36772 71165 36812
rect 73315 36772 73324 36812
rect 73364 36772 73804 36812
rect 73844 36772 73853 36812
rect 73900 36772 76588 36812
rect 76628 36772 77356 36812
rect 77396 36772 77405 36812
rect 0 36728 80 36748
rect 0 36688 38668 36728
rect 38708 36688 38717 36728
rect 57283 36688 57292 36728
rect 57332 36688 58348 36728
rect 58388 36688 58636 36728
rect 58676 36688 58685 36728
rect 60451 36688 60460 36728
rect 60500 36688 61420 36728
rect 61460 36688 63532 36728
rect 63572 36688 63581 36728
rect 63811 36688 63820 36728
rect 63860 36688 64012 36728
rect 64052 36688 64061 36728
rect 65539 36688 65548 36728
rect 65588 36688 66988 36728
rect 67028 36688 67037 36728
rect 68707 36688 68716 36728
rect 68756 36688 69772 36728
rect 69812 36688 69821 36728
rect 72835 36688 72844 36728
rect 72884 36688 75148 36728
rect 75188 36688 76204 36728
rect 76244 36688 76253 36728
rect 76867 36688 76876 36728
rect 76916 36688 78220 36728
rect 78260 36688 78269 36728
rect 0 36668 80 36688
rect 56227 36604 56236 36644
rect 56276 36604 57196 36644
rect 57236 36604 57245 36644
rect 66988 36560 67028 36688
rect 76291 36604 76300 36644
rect 76340 36604 76780 36644
rect 76820 36604 76829 36644
rect 62083 36520 62092 36560
rect 62132 36520 63724 36560
rect 63764 36520 64108 36560
rect 64148 36520 64157 36560
rect 66988 36520 67756 36560
rect 67796 36520 68716 36560
rect 68756 36520 68765 36560
rect 70051 36520 70060 36560
rect 70100 36520 70636 36560
rect 70676 36520 72076 36560
rect 72116 36520 73516 36560
rect 73556 36520 73565 36560
rect 75235 36520 75244 36560
rect 75284 36520 76108 36560
rect 76148 36520 76157 36560
rect 76579 36520 76588 36560
rect 76628 36520 77068 36560
rect 77108 36520 77117 36560
rect 69091 36476 69149 36477
rect 65731 36436 65740 36476
rect 65780 36436 68428 36476
rect 68468 36436 68477 36476
rect 68995 36436 69004 36476
rect 69044 36436 69100 36476
rect 69140 36436 69149 36476
rect 70915 36436 70924 36476
rect 70964 36436 72172 36476
rect 72212 36436 72748 36476
rect 72788 36436 72940 36476
rect 72980 36436 72989 36476
rect 69091 36435 69149 36436
rect 69091 36352 69100 36392
rect 69140 36352 72556 36392
rect 72596 36352 72605 36392
rect 67555 36308 67613 36309
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 15103 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 15489 36308
rect 27103 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 27489 36308
rect 39103 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 39489 36308
rect 51103 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 51489 36308
rect 63103 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 63489 36308
rect 67470 36268 67564 36308
rect 67604 36268 67613 36308
rect 75103 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 75489 36308
rect 67555 36267 67613 36268
rect 76867 36224 76925 36225
rect 67075 36184 67084 36224
rect 67124 36184 69100 36224
rect 69140 36184 69676 36224
rect 69716 36184 69725 36224
rect 74467 36184 74476 36224
rect 74516 36184 76684 36224
rect 76724 36184 76876 36224
rect 76916 36184 76925 36224
rect 76867 36183 76925 36184
rect 69475 36100 69484 36140
rect 69524 36100 70924 36140
rect 70964 36100 70973 36140
rect 71203 36100 71212 36140
rect 71252 36100 71884 36140
rect 71924 36100 74284 36140
rect 74324 36100 74333 36140
rect 76771 36100 76780 36140
rect 76820 36100 77548 36140
rect 77588 36100 77597 36140
rect 49123 36016 49132 36056
rect 49172 36016 50476 36056
rect 50516 36016 50525 36056
rect 61411 36016 61420 36056
rect 61460 36016 62188 36056
rect 62228 36016 62237 36056
rect 68707 36016 68716 36056
rect 68756 36016 70060 36056
rect 70100 36016 70109 36056
rect 73507 36016 73516 36056
rect 73556 36016 74764 36056
rect 74804 36016 75436 36056
rect 75476 36016 78316 36056
rect 78356 36016 78365 36056
rect 43939 35932 43948 35972
rect 43988 35932 50956 35972
rect 50996 35932 56812 35972
rect 56852 35932 56861 35972
rect 60355 35932 60364 35972
rect 60404 35932 61516 35972
rect 61556 35932 61565 35972
rect 66691 35932 66700 35972
rect 66740 35932 68524 35972
rect 68564 35932 68573 35972
rect 73027 35932 73036 35972
rect 73076 35932 73804 35972
rect 73844 35932 75916 35972
rect 75956 35932 75965 35972
rect 0 35828 80 35908
rect 50851 35888 50909 35889
rect 50851 35848 50860 35888
rect 50900 35848 51436 35888
rect 51476 35848 52780 35888
rect 52820 35848 52829 35888
rect 56035 35848 56044 35888
rect 56084 35848 56908 35888
rect 56948 35848 58444 35888
rect 58484 35848 58493 35888
rect 58723 35848 58732 35888
rect 58772 35848 60940 35888
rect 60980 35848 61228 35888
rect 61268 35848 61277 35888
rect 61603 35848 61612 35888
rect 61652 35848 62092 35888
rect 62132 35848 62668 35888
rect 62708 35848 62717 35888
rect 66979 35848 66988 35888
rect 67028 35848 67372 35888
rect 67412 35848 67421 35888
rect 69859 35848 69868 35888
rect 69908 35848 71596 35888
rect 71636 35848 71980 35888
rect 72020 35848 72029 35888
rect 73411 35848 73420 35888
rect 73460 35848 73996 35888
rect 74036 35848 74045 35888
rect 76483 35848 76492 35888
rect 76532 35848 76541 35888
rect 50851 35847 50909 35848
rect 61228 35804 61268 35848
rect 55459 35764 55468 35804
rect 55508 35764 56332 35804
rect 56372 35764 56381 35804
rect 61228 35764 61996 35804
rect 62036 35764 62045 35804
rect 64195 35764 64204 35804
rect 64244 35764 66892 35804
rect 66932 35764 66941 35804
rect 61996 35720 62036 35764
rect 76492 35720 76532 35848
rect 55843 35680 55852 35720
rect 55892 35680 56620 35720
rect 56660 35680 56669 35720
rect 61996 35680 66028 35720
rect 66068 35680 66077 35720
rect 68803 35680 68812 35720
rect 68852 35680 76532 35720
rect 49603 35596 49612 35636
rect 49652 35596 53260 35636
rect 53300 35596 53309 35636
rect 54403 35596 54412 35636
rect 54452 35596 65164 35636
rect 65204 35596 65213 35636
rect 74275 35596 74284 35636
rect 74324 35596 77068 35636
rect 77108 35596 77452 35636
rect 77492 35596 77501 35636
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 16343 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 16729 35552
rect 28343 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 28729 35552
rect 40343 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 40729 35552
rect 52343 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 52729 35552
rect 61411 35512 61420 35552
rect 61460 35512 61708 35552
rect 61748 35512 61757 35552
rect 64343 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 64729 35552
rect 68035 35512 68044 35552
rect 68084 35512 71020 35552
rect 71060 35512 71069 35552
rect 76343 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 76729 35552
rect 70531 35428 70540 35468
rect 70580 35428 70828 35468
rect 70868 35428 73708 35468
rect 73748 35428 78124 35468
rect 78164 35428 78173 35468
rect 55171 35344 55180 35384
rect 55220 35344 55604 35384
rect 65827 35344 65836 35384
rect 65876 35344 66796 35384
rect 66836 35344 66845 35384
rect 77155 35344 77164 35384
rect 77204 35344 77644 35384
rect 77684 35344 77693 35384
rect 55564 35300 55604 35344
rect 51436 35260 51628 35300
rect 51668 35260 54412 35300
rect 54452 35260 54461 35300
rect 54787 35260 54796 35300
rect 54836 35260 55276 35300
rect 55316 35260 55325 35300
rect 55555 35260 55564 35300
rect 55604 35260 55613 35300
rect 66883 35260 66892 35300
rect 66932 35260 67276 35300
rect 67316 35260 67325 35300
rect 70435 35260 70444 35300
rect 70484 35260 71404 35300
rect 71444 35260 71453 35300
rect 72547 35260 72556 35300
rect 72596 35260 73036 35300
rect 73076 35260 73085 35300
rect 51436 35216 51476 35260
rect 51427 35176 51436 35216
rect 51476 35176 51485 35216
rect 52291 35176 52300 35216
rect 52340 35176 55084 35216
rect 55124 35176 55133 35216
rect 56995 35176 57004 35216
rect 57044 35176 58156 35216
rect 58196 35176 58205 35216
rect 66115 35176 66124 35216
rect 66164 35176 66604 35216
rect 66644 35176 66796 35216
rect 66836 35176 66845 35216
rect 68227 35176 68236 35216
rect 68276 35176 70540 35216
rect 70580 35176 70589 35216
rect 70723 35176 70732 35216
rect 70772 35176 71884 35216
rect 71924 35176 71933 35216
rect 72739 35176 72748 35216
rect 72788 35176 72797 35216
rect 74179 35176 74188 35216
rect 74228 35176 76108 35216
rect 76148 35176 76157 35216
rect 77443 35176 77452 35216
rect 77492 35176 77836 35216
rect 77876 35176 77885 35216
rect 72748 35132 72788 35176
rect 51523 35092 51532 35132
rect 51572 35092 52108 35132
rect 52148 35092 52157 35132
rect 55843 35092 55852 35132
rect 55892 35092 56044 35132
rect 56084 35092 56093 35132
rect 72748 35092 73228 35132
rect 73268 35092 73460 35132
rect 0 34988 80 35068
rect 73420 35048 73460 35092
rect 50467 35008 50476 35048
rect 50516 35008 51340 35048
rect 51380 35008 51389 35048
rect 61411 35008 61420 35048
rect 61460 35008 65932 35048
rect 65972 35008 65981 35048
rect 71683 35008 71692 35048
rect 71732 35008 72364 35048
rect 72404 35008 72413 35048
rect 72547 35008 72556 35048
rect 72596 35008 72748 35048
rect 72788 35008 72797 35048
rect 73420 35008 76492 35048
rect 76532 35008 76876 35048
rect 76916 35008 76925 35048
rect 57475 34924 57484 34964
rect 57524 34924 58156 34964
rect 58196 34924 58205 34964
rect 72067 34924 72076 34964
rect 72116 34924 72460 34964
rect 72500 34924 72509 34964
rect 56419 34840 56428 34880
rect 56468 34840 57964 34880
rect 58004 34840 69196 34880
rect 69236 34840 69245 34880
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 15103 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 15489 34796
rect 27103 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 27489 34796
rect 39103 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 39489 34796
rect 51103 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 51489 34796
rect 55171 34756 55180 34796
rect 55220 34756 58196 34796
rect 62179 34756 62188 34796
rect 62228 34756 62668 34796
rect 62708 34756 62717 34796
rect 63103 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 63489 34796
rect 75103 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 75489 34796
rect 50371 34672 50380 34712
rect 50420 34672 51724 34712
rect 51764 34672 51773 34712
rect 52771 34672 52780 34712
rect 52820 34672 54988 34712
rect 55028 34672 55037 34712
rect 58156 34628 58196 34756
rect 61507 34672 61516 34712
rect 61556 34672 64108 34712
rect 64148 34672 64157 34712
rect 66979 34672 66988 34712
rect 67028 34672 67468 34712
rect 67508 34672 67517 34712
rect 51139 34588 51148 34628
rect 51188 34588 51532 34628
rect 51572 34588 51581 34628
rect 58147 34588 58156 34628
rect 58196 34588 59116 34628
rect 59156 34588 59165 34628
rect 66691 34588 66700 34628
rect 66740 34588 67660 34628
rect 67700 34588 67709 34628
rect 68899 34588 68908 34628
rect 68948 34588 69964 34628
rect 70004 34588 70444 34628
rect 70484 34588 70493 34628
rect 77932 34588 78124 34628
rect 78164 34588 78173 34628
rect 45955 34504 45964 34544
rect 46004 34504 46540 34544
rect 46580 34504 46589 34544
rect 46819 34504 46828 34544
rect 46868 34504 49228 34544
rect 49268 34504 49277 34544
rect 51235 34504 51244 34544
rect 51284 34504 52204 34544
rect 52244 34504 52253 34544
rect 55939 34504 55948 34544
rect 55988 34504 56524 34544
rect 56564 34504 56573 34544
rect 58339 34504 58348 34544
rect 58388 34504 58397 34544
rect 59779 34504 59788 34544
rect 59828 34504 61900 34544
rect 61940 34504 61949 34544
rect 62563 34504 62572 34544
rect 62612 34504 63380 34544
rect 66403 34504 66412 34544
rect 66452 34504 66740 34544
rect 68035 34504 68044 34544
rect 68084 34504 70348 34544
rect 70388 34504 70636 34544
rect 70676 34504 70685 34544
rect 71299 34504 71308 34544
rect 71348 34504 71788 34544
rect 71828 34504 71837 34544
rect 55948 34420 56428 34460
rect 56468 34420 56477 34460
rect 55948 34376 55988 34420
rect 48451 34336 48460 34376
rect 48500 34336 49516 34376
rect 49556 34336 50476 34376
rect 50516 34336 50525 34376
rect 51811 34336 51820 34376
rect 51860 34336 52396 34376
rect 52436 34336 52445 34376
rect 54115 34336 54124 34376
rect 54164 34336 55084 34376
rect 55124 34336 55133 34376
rect 55939 34336 55948 34376
rect 55988 34336 55997 34376
rect 56227 34336 56236 34376
rect 56276 34336 58252 34376
rect 58292 34336 58301 34376
rect 58348 34292 58388 34504
rect 63340 34460 63380 34504
rect 66700 34460 66740 34504
rect 59587 34420 59596 34460
rect 59636 34420 60172 34460
rect 60212 34420 60221 34460
rect 62659 34420 62668 34460
rect 62708 34420 63244 34460
rect 63284 34420 63293 34460
rect 63340 34420 63628 34460
rect 63668 34420 63677 34460
rect 66691 34420 66700 34460
rect 66740 34420 66749 34460
rect 68995 34420 69004 34460
rect 69044 34420 72020 34460
rect 71980 34376 72020 34420
rect 77932 34376 77972 34588
rect 59203 34336 59212 34376
rect 59252 34336 59980 34376
rect 60020 34336 61036 34376
rect 61076 34336 61085 34376
rect 62083 34336 62092 34376
rect 62132 34336 62764 34376
rect 62804 34336 62813 34376
rect 67267 34336 67276 34376
rect 67316 34336 67564 34376
rect 67604 34336 67613 34376
rect 67660 34336 67669 34376
rect 67709 34336 69868 34376
rect 69908 34336 69917 34376
rect 71971 34336 71980 34376
rect 72020 34336 72029 34376
rect 76195 34336 76204 34376
rect 76244 34336 77644 34376
rect 77684 34336 77693 34376
rect 77923 34336 77932 34376
rect 77972 34336 77981 34376
rect 78115 34336 78124 34376
rect 78164 34336 79468 34376
rect 79508 34336 79517 34376
rect 78124 34292 78164 34336
rect 56323 34252 56332 34292
rect 56372 34252 58828 34292
rect 58868 34252 58877 34292
rect 62659 34252 62668 34292
rect 62708 34252 63052 34292
rect 63092 34252 63101 34292
rect 67459 34252 67468 34292
rect 67508 34252 67517 34292
rect 76867 34252 76876 34292
rect 76916 34252 77356 34292
rect 77396 34252 78164 34292
rect 0 34148 80 34228
rect 67468 34208 67508 34252
rect 52483 34168 52492 34208
rect 52532 34168 53644 34208
rect 53684 34168 53693 34208
rect 58051 34168 58060 34208
rect 58100 34168 58444 34208
rect 58484 34168 58493 34208
rect 66211 34168 66220 34208
rect 66260 34168 66796 34208
rect 66836 34168 66845 34208
rect 67171 34168 67180 34208
rect 67220 34168 67508 34208
rect 71395 34168 71404 34208
rect 71444 34168 71788 34208
rect 71828 34168 74572 34208
rect 74612 34168 75628 34208
rect 75668 34168 75677 34208
rect 49219 34084 49228 34124
rect 49268 34084 50092 34124
rect 50132 34084 52204 34124
rect 52244 34084 54124 34124
rect 54164 34084 54173 34124
rect 63235 34084 63244 34124
rect 63284 34084 65452 34124
rect 65492 34084 69580 34124
rect 69620 34084 69629 34124
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 16343 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 16729 34040
rect 28343 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 28729 34040
rect 40343 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 40729 34040
rect 52343 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 52729 34040
rect 55843 34000 55852 34040
rect 55892 34000 56236 34040
rect 56276 34000 56285 34040
rect 62083 34000 62092 34040
rect 62132 34000 62572 34040
rect 62612 34000 62621 34040
rect 62851 34000 62860 34040
rect 62900 34000 63148 34040
rect 63188 34000 63197 34040
rect 64343 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 64729 34040
rect 76343 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 76729 34040
rect 67555 33956 67613 33957
rect 54595 33916 54604 33956
rect 54644 33916 55276 33956
rect 55316 33916 55325 33956
rect 57763 33916 57772 33956
rect 57812 33916 58348 33956
rect 58388 33916 58397 33956
rect 63052 33916 66316 33956
rect 66356 33916 67180 33956
rect 67220 33916 67229 33956
rect 67470 33916 67564 33956
rect 67604 33916 67613 33956
rect 69859 33916 69868 33956
rect 69908 33916 73708 33956
rect 73748 33916 73757 33956
rect 55075 33832 55084 33872
rect 55124 33832 55316 33872
rect 52195 33748 52204 33788
rect 52244 33748 54028 33788
rect 54068 33748 54077 33788
rect 49123 33664 49132 33704
rect 49172 33664 50956 33704
rect 50996 33664 51005 33704
rect 53635 33580 53644 33620
rect 53684 33580 54604 33620
rect 54644 33580 54653 33620
rect 55276 33536 55316 33832
rect 63052 33788 63092 33916
rect 67555 33915 67613 33916
rect 71971 33832 71980 33872
rect 72020 33832 77260 33872
rect 77300 33832 77309 33872
rect 76867 33788 76925 33789
rect 57571 33748 57580 33788
rect 57620 33748 57772 33788
rect 57812 33748 57821 33788
rect 60163 33748 60172 33788
rect 60212 33748 63052 33788
rect 63092 33748 63101 33788
rect 76782 33748 76876 33788
rect 76916 33748 76925 33788
rect 76867 33747 76925 33748
rect 59683 33664 59692 33704
rect 59732 33664 61612 33704
rect 61652 33664 62380 33704
rect 62420 33664 62429 33704
rect 71587 33664 71596 33704
rect 71636 33664 72460 33704
rect 72500 33664 72509 33704
rect 74851 33664 74860 33704
rect 74900 33664 76300 33704
rect 76340 33664 76349 33704
rect 76483 33664 76492 33704
rect 76532 33664 76972 33704
rect 77012 33664 77021 33704
rect 77443 33664 77452 33704
rect 77492 33664 78412 33704
rect 78452 33664 78461 33704
rect 77452 33620 77492 33664
rect 61315 33580 61324 33620
rect 61364 33580 62188 33620
rect 62228 33580 66124 33620
rect 66164 33580 66173 33620
rect 72259 33580 72268 33620
rect 72308 33580 72556 33620
rect 72596 33580 72605 33620
rect 75811 33580 75820 33620
rect 75860 33580 77492 33620
rect 55267 33496 55276 33536
rect 55316 33496 55325 33536
rect 61123 33496 61132 33536
rect 61172 33496 62476 33536
rect 62516 33496 62525 33536
rect 65923 33496 65932 33536
rect 65972 33496 66220 33536
rect 66260 33496 66269 33536
rect 75523 33496 75532 33536
rect 75572 33496 76396 33536
rect 76436 33496 76445 33536
rect 51523 33412 51532 33452
rect 51572 33412 51820 33452
rect 51860 33412 54796 33452
rect 54836 33412 54845 33452
rect 58531 33412 58540 33452
rect 58580 33412 58924 33452
rect 58964 33412 58973 33452
rect 74755 33412 74764 33452
rect 74804 33412 76012 33452
rect 76052 33412 76061 33452
rect 76771 33412 76780 33452
rect 76820 33412 77548 33452
rect 77588 33412 77597 33452
rect 0 33308 80 33388
rect 54883 33328 54892 33368
rect 54932 33328 55372 33368
rect 55412 33328 55421 33368
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 15103 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 15489 33284
rect 27103 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 27489 33284
rect 39103 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 39489 33284
rect 43171 33244 43180 33284
rect 43220 33244 43948 33284
rect 43988 33244 43997 33284
rect 51103 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 51489 33284
rect 54307 33244 54316 33284
rect 54356 33244 56332 33284
rect 56372 33244 56381 33284
rect 58723 33244 58732 33284
rect 58772 33244 60364 33284
rect 60404 33244 60413 33284
rect 63103 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 63489 33284
rect 75103 33244 75112 33284
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75480 33244 75489 33284
rect 43180 33200 43220 33244
rect 42115 33160 42124 33200
rect 42164 33160 43220 33200
rect 46723 33160 46732 33200
rect 46772 33160 48556 33200
rect 48596 33160 48605 33200
rect 55651 33160 55660 33200
rect 55700 33160 55740 33200
rect 70339 33160 70348 33200
rect 70388 33160 74860 33200
rect 74900 33160 74909 33200
rect 55660 33116 55700 33160
rect 45859 33076 45868 33116
rect 45908 33076 46828 33116
rect 46868 33076 47596 33116
rect 47636 33076 47645 33116
rect 49027 33076 49036 33116
rect 49076 33076 50572 33116
rect 50612 33076 53740 33116
rect 53780 33076 53789 33116
rect 54595 33076 54604 33116
rect 54644 33076 55700 33116
rect 59107 33076 59116 33116
rect 59156 33076 59404 33116
rect 59444 33076 62860 33116
rect 62900 33076 64108 33116
rect 64148 33076 64157 33116
rect 61516 33032 61556 33076
rect 48067 32992 48076 33032
rect 48116 32992 48652 33032
rect 48692 32992 48701 33032
rect 48931 32992 48940 33032
rect 48980 32992 50092 33032
rect 50132 32992 50668 33032
rect 50708 32992 51148 33032
rect 51188 32992 51197 33032
rect 53260 32992 57676 33032
rect 57716 32992 57725 33032
rect 60739 32992 60748 33032
rect 60788 32992 61324 33032
rect 61364 32992 61373 33032
rect 61507 32992 61516 33032
rect 61556 32992 61596 33032
rect 53260 32948 53300 32992
rect 42211 32908 42220 32948
rect 42260 32908 42796 32948
rect 42836 32908 53300 32948
rect 62467 32908 62476 32948
rect 62516 32908 64012 32948
rect 64052 32908 64061 32948
rect 71107 32908 71116 32948
rect 71156 32908 73132 32948
rect 73172 32908 73181 32948
rect 50851 32864 50909 32865
rect 46915 32824 46924 32864
rect 46964 32824 47692 32864
rect 47732 32824 47741 32864
rect 48259 32824 48268 32864
rect 48308 32824 48844 32864
rect 48884 32824 48893 32864
rect 50766 32824 50860 32864
rect 50900 32824 50909 32864
rect 51139 32824 51148 32864
rect 51188 32824 53836 32864
rect 53876 32824 53885 32864
rect 54883 32824 54892 32864
rect 54932 32824 55180 32864
rect 55220 32824 55229 32864
rect 57763 32824 57772 32864
rect 57812 32824 58444 32864
rect 58484 32824 58493 32864
rect 62275 32824 62284 32864
rect 62324 32824 62572 32864
rect 62612 32824 62621 32864
rect 66019 32824 66028 32864
rect 66068 32824 68620 32864
rect 68660 32824 68812 32864
rect 68852 32824 68861 32864
rect 72547 32824 72556 32864
rect 72596 32824 72844 32864
rect 72884 32824 72893 32864
rect 77155 32824 77164 32864
rect 77204 32824 77836 32864
rect 77876 32824 77885 32864
rect 78115 32824 78124 32864
rect 78164 32824 78508 32864
rect 78548 32824 78557 32864
rect 50851 32823 50909 32824
rect 50860 32780 50900 32823
rect 45955 32740 45964 32780
rect 46004 32740 47212 32780
rect 47252 32740 47261 32780
rect 50860 32740 51820 32780
rect 51860 32740 51869 32780
rect 58339 32740 58348 32780
rect 58388 32740 58732 32780
rect 58772 32740 58781 32780
rect 50563 32656 50572 32696
rect 50612 32656 51244 32696
rect 51284 32656 51293 32696
rect 65635 32656 65644 32696
rect 65684 32656 66260 32696
rect 68995 32656 69004 32696
rect 69044 32656 69772 32696
rect 69812 32656 69821 32696
rect 70531 32656 70540 32696
rect 70580 32656 70828 32696
rect 70868 32656 71692 32696
rect 71732 32656 71980 32696
rect 72020 32656 72029 32696
rect 75820 32656 76588 32696
rect 76628 32656 76637 32696
rect 66220 32612 66260 32656
rect 70627 32612 70685 32613
rect 54979 32572 54988 32612
rect 55028 32572 58060 32612
rect 58100 32572 65932 32612
rect 65972 32572 65981 32612
rect 66220 32572 70636 32612
rect 70676 32572 70685 32612
rect 70627 32571 70685 32572
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 16343 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 16729 32528
rect 28343 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 28729 32528
rect 40343 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 40729 32528
rect 52343 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 52729 32528
rect 54691 32488 54700 32528
rect 54740 32488 55564 32528
rect 55604 32488 55613 32528
rect 58627 32488 58636 32528
rect 58676 32488 59020 32528
rect 59060 32488 59069 32528
rect 62659 32488 62668 32528
rect 62708 32488 63436 32528
rect 63476 32488 63485 32528
rect 64343 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 64729 32528
rect 65347 32488 65356 32528
rect 65396 32488 66892 32528
rect 66932 32488 66941 32528
rect 69091 32488 69100 32528
rect 69140 32488 69676 32528
rect 69716 32488 71116 32528
rect 71156 32488 71165 32528
rect 72067 32488 72076 32528
rect 72116 32488 72940 32528
rect 72980 32488 72989 32528
rect 46531 32404 46540 32444
rect 46580 32404 47308 32444
rect 47348 32404 48268 32444
rect 48308 32404 66220 32444
rect 66260 32404 66269 32444
rect 68899 32404 68908 32444
rect 68948 32404 70924 32444
rect 70964 32404 71500 32444
rect 71540 32404 71549 32444
rect 46243 32320 46252 32360
rect 46292 32320 46636 32360
rect 46676 32320 46685 32360
rect 58819 32320 58828 32360
rect 58868 32320 59596 32360
rect 59636 32320 59645 32360
rect 63340 32320 64492 32360
rect 64532 32320 65644 32360
rect 65684 32320 65693 32360
rect 66883 32320 66892 32360
rect 66932 32320 67180 32360
rect 67220 32320 67229 32360
rect 69283 32320 69292 32360
rect 69332 32320 69964 32360
rect 70004 32320 70013 32360
rect 71011 32320 71020 32360
rect 71060 32320 71596 32360
rect 71636 32320 71645 32360
rect 71875 32320 71884 32360
rect 71924 32320 72652 32360
rect 72692 32320 72940 32360
rect 72980 32320 72989 32360
rect 63340 32276 63380 32320
rect 58339 32236 58348 32276
rect 58388 32236 63052 32276
rect 63092 32236 63101 32276
rect 63235 32236 63244 32276
rect 63284 32236 63380 32276
rect 64099 32236 64108 32276
rect 64148 32236 64780 32276
rect 64820 32236 65356 32276
rect 65396 32236 65405 32276
rect 71107 32236 71116 32276
rect 71156 32236 73460 32276
rect 73420 32192 73460 32236
rect 75820 32192 75860 32656
rect 76343 32488 76352 32528
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76720 32488 76729 32528
rect 76003 32320 76012 32360
rect 76052 32320 76300 32360
rect 76340 32320 76349 32360
rect 76483 32320 76492 32360
rect 76532 32320 77452 32360
rect 77492 32320 77501 32360
rect 76867 32276 76925 32277
rect 76012 32236 76684 32276
rect 76724 32236 76876 32276
rect 76916 32236 76925 32276
rect 76012 32192 76052 32236
rect 76867 32235 76925 32236
rect 77443 32192 77501 32193
rect 47107 32152 47116 32192
rect 47156 32152 47404 32192
rect 47444 32152 48460 32192
rect 48500 32152 49612 32192
rect 49652 32152 49661 32192
rect 52387 32152 52396 32192
rect 52436 32152 53452 32192
rect 53492 32152 53501 32192
rect 54220 32152 72748 32192
rect 72788 32152 72797 32192
rect 73420 32152 75820 32192
rect 75860 32152 75869 32192
rect 76003 32152 76012 32192
rect 76052 32152 76061 32192
rect 76867 32152 76876 32192
rect 76916 32152 77452 32192
rect 77492 32152 77740 32192
rect 77780 32152 79468 32192
rect 79508 32152 79517 32192
rect 54220 32108 54260 32152
rect 77443 32151 77501 32152
rect 45667 32068 45676 32108
rect 45716 32068 46540 32108
rect 46580 32068 46589 32108
rect 49123 32068 49132 32108
rect 49172 32068 49420 32108
rect 49460 32068 54260 32108
rect 54403 32068 54412 32108
rect 54452 32068 54892 32108
rect 54932 32068 55180 32108
rect 55220 32068 55229 32108
rect 58435 32068 58444 32108
rect 58484 32068 59308 32108
rect 59348 32068 59357 32108
rect 61603 32068 61612 32108
rect 61652 32068 61900 32108
rect 61940 32068 61949 32108
rect 62467 32068 62476 32108
rect 62516 32068 64340 32108
rect 72643 32068 72652 32108
rect 72692 32068 73036 32108
rect 73076 32068 73085 32108
rect 64300 32024 64340 32068
rect 42499 31984 42508 32024
rect 42548 31984 42644 32024
rect 50563 31984 50572 32024
rect 50612 31984 53548 32024
rect 53588 31984 64244 32024
rect 64291 31984 64300 32024
rect 64340 31984 64349 32024
rect 65443 31984 65452 32024
rect 65492 31984 66604 32024
rect 66644 31984 66653 32024
rect 69859 31984 69868 32024
rect 69908 31984 72172 32024
rect 72212 31984 72556 32024
rect 72596 31984 72605 32024
rect 42604 31772 42644 31984
rect 64204 31940 64244 31984
rect 54787 31900 54796 31940
rect 54836 31900 55756 31940
rect 55796 31900 55805 31940
rect 62851 31900 62860 31940
rect 62900 31900 63532 31940
rect 63572 31900 64012 31940
rect 64052 31900 64061 31940
rect 64204 31900 65164 31940
rect 65204 31900 65213 31940
rect 66115 31900 66124 31940
rect 66164 31900 67084 31940
rect 67124 31900 67133 31940
rect 49027 31816 49036 31856
rect 49076 31816 50036 31856
rect 58627 31816 58636 31856
rect 58676 31816 61132 31856
rect 61172 31816 67852 31856
rect 67892 31816 67901 31856
rect 72931 31816 72940 31856
rect 72980 31816 74572 31856
rect 74612 31816 74621 31856
rect 49996 31772 50036 31816
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 15103 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 15489 31772
rect 27103 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 27489 31772
rect 39103 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 39489 31772
rect 41740 31732 42644 31772
rect 48835 31732 48844 31772
rect 48884 31732 49228 31772
rect 49268 31732 49277 31772
rect 49987 31732 49996 31772
rect 50036 31732 50668 31772
rect 50708 31732 50717 31772
rect 51103 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 51489 31772
rect 59107 31732 59116 31772
rect 59156 31732 60460 31772
rect 60500 31732 60509 31772
rect 63103 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 63489 31772
rect 72355 31732 72364 31772
rect 72404 31732 74284 31772
rect 74324 31732 74333 31772
rect 75103 31732 75112 31772
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75480 31732 75489 31772
rect 0 31628 80 31708
rect 41740 31688 41780 31732
rect 42604 31688 42644 31732
rect 40963 31648 40972 31688
rect 41012 31648 41780 31688
rect 41827 31648 41836 31688
rect 41876 31648 42508 31688
rect 42548 31648 42557 31688
rect 42604 31648 45004 31688
rect 45044 31648 45053 31688
rect 59011 31648 59020 31688
rect 59060 31648 59980 31688
rect 60020 31648 61900 31688
rect 61940 31648 64204 31688
rect 64244 31648 64253 31688
rect 69475 31648 69484 31688
rect 69524 31648 70636 31688
rect 70676 31648 73036 31688
rect 73076 31648 73324 31688
rect 73364 31648 73373 31688
rect 74851 31648 74860 31688
rect 74900 31648 76204 31688
rect 76244 31648 78316 31688
rect 78356 31648 78365 31688
rect 42307 31564 42316 31604
rect 42356 31564 43084 31604
rect 43124 31564 46060 31604
rect 46100 31564 46109 31604
rect 59683 31564 59692 31604
rect 59732 31564 60076 31604
rect 60116 31564 60125 31604
rect 70723 31564 70732 31604
rect 70772 31564 71116 31604
rect 71156 31564 71165 31604
rect 49507 31480 49516 31520
rect 49556 31480 49708 31520
rect 49748 31480 49757 31520
rect 59779 31480 59788 31520
rect 59828 31480 59980 31520
rect 60020 31480 60029 31520
rect 68611 31480 68620 31520
rect 68660 31480 68812 31520
rect 68852 31480 68861 31520
rect 76195 31480 76204 31520
rect 76244 31480 76492 31520
rect 76532 31480 76541 31520
rect 51619 31436 51677 31437
rect 71971 31436 72029 31437
rect 42979 31396 42988 31436
rect 43028 31396 43220 31436
rect 51534 31396 51628 31436
rect 51668 31396 51677 31436
rect 51907 31396 51916 31436
rect 51956 31396 55468 31436
rect 55508 31396 55517 31436
rect 63349 31396 63358 31436
rect 63398 31396 64396 31436
rect 64436 31396 64445 31436
rect 66403 31396 66412 31436
rect 66452 31396 66796 31436
rect 66836 31396 66988 31436
rect 67028 31396 67037 31436
rect 70915 31396 70924 31436
rect 70964 31396 71980 31436
rect 72020 31396 72029 31436
rect 43180 31352 43220 31396
rect 51619 31395 51677 31396
rect 71971 31395 72029 31396
rect 43180 31312 43756 31352
rect 43796 31312 43805 31352
rect 46147 31312 46156 31352
rect 46196 31312 47212 31352
rect 47252 31312 48652 31352
rect 48692 31312 49324 31352
rect 49364 31312 49373 31352
rect 51139 31312 51148 31352
rect 51188 31312 52108 31352
rect 52148 31312 52157 31352
rect 53443 31312 53452 31352
rect 53492 31312 54028 31352
rect 54068 31312 56908 31352
rect 56948 31312 57388 31352
rect 57428 31312 59020 31352
rect 59060 31312 59069 31352
rect 60451 31312 60460 31352
rect 60500 31312 62092 31352
rect 62132 31312 63052 31352
rect 63092 31312 63101 31352
rect 70723 31312 70732 31352
rect 70772 31312 71308 31352
rect 71348 31312 71357 31352
rect 73027 31312 73036 31352
rect 73076 31312 74668 31352
rect 74708 31312 74717 31352
rect 76771 31312 76780 31352
rect 76820 31312 77164 31352
rect 77204 31312 78220 31352
rect 78260 31312 78269 31352
rect 77251 31268 77309 31269
rect 60355 31228 60364 31268
rect 60404 31228 62668 31268
rect 62708 31228 62717 31268
rect 66691 31228 66700 31268
rect 66740 31228 66988 31268
rect 67028 31228 67037 31268
rect 77059 31228 77068 31268
rect 77108 31228 77260 31268
rect 77300 31228 77309 31268
rect 77251 31227 77309 31228
rect 71107 31184 71165 31185
rect 76867 31184 76925 31185
rect 41923 31144 41932 31184
rect 41972 31144 42508 31184
rect 42548 31144 42988 31184
rect 43028 31144 43037 31184
rect 48067 31144 48076 31184
rect 48116 31144 49324 31184
rect 49364 31144 49373 31184
rect 70435 31144 70444 31184
rect 70484 31144 70828 31184
rect 70868 31144 70877 31184
rect 71022 31144 71116 31184
rect 71156 31144 71165 31184
rect 76099 31144 76108 31184
rect 76148 31144 76300 31184
rect 76340 31144 76349 31184
rect 76867 31144 76876 31184
rect 76916 31144 77452 31184
rect 77492 31144 77501 31184
rect 71107 31143 71165 31144
rect 76867 31143 76925 31144
rect 77164 31100 77204 31144
rect 56611 31060 56620 31100
rect 56660 31060 58540 31100
rect 58580 31060 66604 31100
rect 66644 31060 66653 31100
rect 67075 31060 67084 31100
rect 67124 31060 69100 31100
rect 69140 31060 73516 31100
rect 73556 31060 73565 31100
rect 77155 31060 77164 31100
rect 77204 31060 77244 31100
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 16343 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 16729 31016
rect 28343 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 28729 31016
rect 40343 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 40729 31016
rect 43363 30976 43372 31016
rect 43412 30976 43421 31016
rect 43939 30976 43948 31016
rect 43988 30976 48844 31016
rect 48884 30976 48893 31016
rect 52343 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 52729 31016
rect 55267 30976 55276 31016
rect 55316 30976 55948 31016
rect 55988 30976 55997 31016
rect 64343 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 64729 31016
rect 76343 30976 76352 31016
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76720 30976 76729 31016
rect 43372 30932 43412 30976
rect 42019 30892 42028 30932
rect 42068 30892 43412 30932
rect 45091 30892 45100 30932
rect 45140 30892 46348 30932
rect 46388 30892 46397 30932
rect 0 30788 80 30868
rect 43180 30848 43220 30892
rect 42211 30808 42220 30848
rect 42260 30808 42508 30848
rect 42548 30808 42557 30848
rect 43180 30808 47636 30848
rect 49411 30808 49420 30848
rect 49460 30808 50860 30848
rect 50900 30808 50909 30848
rect 52099 30808 52108 30848
rect 52148 30808 55948 30848
rect 55988 30808 58156 30848
rect 58196 30808 58205 30848
rect 70540 30808 71212 30848
rect 71252 30808 71261 30848
rect 73603 30808 73612 30848
rect 73652 30808 75436 30848
rect 75476 30808 75485 30848
rect 44995 30724 45004 30764
rect 45044 30724 46444 30764
rect 46484 30724 46493 30764
rect 44227 30640 44236 30680
rect 44276 30640 44908 30680
rect 44948 30640 44957 30680
rect 46051 30640 46060 30680
rect 46100 30640 47500 30680
rect 47540 30640 47549 30680
rect 41155 30596 41213 30597
rect 47596 30596 47636 30808
rect 49891 30724 49900 30764
rect 49940 30724 50380 30764
rect 50420 30724 51148 30764
rect 51188 30724 51724 30764
rect 51764 30724 51773 30764
rect 55363 30724 55372 30764
rect 55412 30724 56620 30764
rect 56660 30724 56669 30764
rect 57763 30724 57772 30764
rect 57812 30724 59692 30764
rect 59732 30724 59741 30764
rect 65827 30724 65836 30764
rect 65876 30724 66124 30764
rect 66164 30724 66173 30764
rect 70540 30680 70580 30808
rect 70627 30724 70636 30764
rect 70676 30724 71308 30764
rect 71348 30724 71357 30764
rect 74851 30724 74860 30764
rect 74900 30724 75340 30764
rect 75380 30724 75389 30764
rect 76483 30724 76492 30764
rect 76532 30724 77644 30764
rect 77684 30724 77693 30764
rect 50755 30640 50764 30680
rect 50804 30640 51820 30680
rect 51860 30640 51869 30680
rect 54691 30640 54700 30680
rect 54740 30640 55660 30680
rect 55700 30640 56140 30680
rect 56180 30640 56189 30680
rect 59692 30640 60076 30680
rect 60116 30640 61132 30680
rect 61172 30640 62476 30680
rect 62516 30640 62860 30680
rect 62900 30640 62909 30680
rect 63715 30640 63724 30680
rect 63764 30640 63956 30680
rect 64387 30640 64396 30680
rect 64436 30640 67276 30680
rect 67316 30640 67948 30680
rect 67988 30640 68908 30680
rect 68948 30640 69484 30680
rect 69524 30640 69533 30680
rect 70531 30640 70540 30680
rect 70580 30640 70589 30680
rect 75139 30640 75148 30680
rect 75188 30640 76012 30680
rect 76052 30640 76588 30680
rect 76628 30640 76637 30680
rect 77443 30640 77452 30680
rect 77492 30640 77836 30680
rect 77876 30640 77885 30680
rect 59692 30596 59732 30640
rect 63916 30596 63956 30640
rect 71971 30596 72029 30597
rect 77251 30596 77309 30597
rect 3811 30556 3820 30596
rect 3860 30556 40588 30596
rect 40628 30556 40637 30596
rect 41070 30556 41164 30596
rect 41204 30556 41213 30596
rect 42115 30556 42124 30596
rect 42164 30556 42412 30596
rect 42452 30556 42461 30596
rect 43267 30556 43276 30596
rect 43316 30556 45676 30596
rect 45716 30556 45725 30596
rect 46531 30556 46540 30596
rect 46580 30556 47116 30596
rect 47156 30556 47165 30596
rect 47596 30556 51532 30596
rect 51572 30556 52204 30596
rect 52244 30556 52253 30596
rect 56227 30556 56236 30596
rect 56276 30556 56524 30596
rect 56564 30556 56573 30596
rect 59683 30556 59692 30596
rect 59732 30556 59741 30596
rect 60739 30556 60748 30596
rect 60788 30556 62284 30596
rect 62324 30556 63820 30596
rect 63860 30556 63869 30596
rect 63916 30556 64204 30596
rect 64244 30556 65932 30596
rect 65972 30556 71980 30596
rect 72020 30556 72029 30596
rect 75523 30556 75532 30596
rect 75572 30556 77260 30596
rect 77300 30556 77309 30596
rect 41155 30555 41213 30556
rect 71971 30555 72029 30556
rect 77251 30555 77309 30556
rect 43075 30472 43084 30512
rect 43124 30472 43948 30512
rect 43988 30472 43997 30512
rect 48835 30472 48844 30512
rect 48884 30472 49420 30512
rect 49460 30472 49469 30512
rect 51619 30472 51628 30512
rect 51668 30472 52300 30512
rect 52340 30472 52349 30512
rect 52771 30472 52780 30512
rect 52820 30472 54508 30512
rect 54548 30472 54557 30512
rect 71395 30472 71404 30512
rect 71444 30472 72652 30512
rect 72692 30472 76492 30512
rect 76532 30472 76780 30512
rect 76820 30472 76829 30512
rect 77635 30472 77644 30512
rect 77684 30472 77836 30512
rect 77876 30472 79468 30512
rect 79508 30472 79517 30512
rect 40099 30388 40108 30428
rect 40148 30388 42796 30428
rect 42836 30388 42845 30428
rect 45283 30388 45292 30428
rect 45332 30388 45964 30428
rect 46004 30388 46348 30428
rect 46388 30388 46397 30428
rect 50755 30388 50764 30428
rect 50804 30388 51244 30428
rect 51284 30388 51293 30428
rect 51715 30388 51724 30428
rect 51764 30388 55084 30428
rect 55124 30388 55133 30428
rect 60931 30388 60940 30428
rect 60980 30388 61076 30428
rect 71203 30388 71212 30428
rect 71252 30388 72172 30428
rect 72212 30388 73708 30428
rect 73748 30388 74188 30428
rect 74228 30388 74237 30428
rect 51724 30344 51764 30388
rect 40972 30304 41836 30344
rect 41876 30304 42604 30344
rect 42644 30304 45100 30344
rect 45140 30304 45149 30344
rect 50275 30304 50284 30344
rect 50324 30304 51764 30344
rect 55939 30304 55948 30344
rect 55988 30304 56332 30344
rect 56372 30304 56381 30344
rect 40972 30260 41012 30304
rect 61036 30260 61076 30388
rect 72451 30260 72509 30261
rect 76099 30260 76157 30261
rect 77251 30260 77309 30261
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 15103 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 15489 30260
rect 27103 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 27489 30260
rect 39103 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 39489 30260
rect 40963 30220 40972 30260
rect 41012 30220 41021 30260
rect 41347 30220 41356 30260
rect 41396 30220 44524 30260
rect 44564 30220 44573 30260
rect 49315 30220 49324 30260
rect 49364 30220 49373 30260
rect 51103 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 51489 30260
rect 51715 30220 51724 30260
rect 51764 30220 52108 30260
rect 52148 30220 52157 30260
rect 54979 30220 54988 30260
rect 55028 30220 56236 30260
rect 56276 30220 56285 30260
rect 59779 30220 59788 30260
rect 59828 30220 60940 30260
rect 60980 30220 60989 30260
rect 61036 30220 61268 30260
rect 63103 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 63489 30260
rect 63532 30220 65356 30260
rect 65396 30220 65548 30260
rect 65588 30220 65597 30260
rect 71683 30220 71692 30260
rect 71732 30220 71741 30260
rect 72366 30220 72460 30260
rect 72500 30220 72509 30260
rect 75103 30220 75112 30260
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75480 30220 75489 30260
rect 76014 30220 76108 30260
rect 76148 30220 76157 30260
rect 77166 30220 77260 30260
rect 77300 30220 77309 30260
rect 49324 30176 49364 30220
rect 39532 30136 40588 30176
rect 40628 30136 41836 30176
rect 41876 30136 44140 30176
rect 44180 30136 46156 30176
rect 46196 30136 46205 30176
rect 47779 30136 47788 30176
rect 47828 30136 52492 30176
rect 52532 30136 52541 30176
rect 60547 30136 60556 30176
rect 60596 30136 61132 30176
rect 61172 30136 61181 30176
rect 39532 30092 39572 30136
rect 40771 30092 40829 30093
rect 39523 30052 39532 30092
rect 39572 30052 39581 30092
rect 40771 30052 40780 30092
rect 40820 30052 41644 30092
rect 41684 30052 44044 30092
rect 44084 30052 44093 30092
rect 44899 30052 44908 30092
rect 44948 30052 45964 30092
rect 46004 30052 46013 30092
rect 58339 30052 58348 30092
rect 58388 30052 58828 30092
rect 58868 30052 58877 30092
rect 59299 30052 59308 30092
rect 59348 30052 59357 30092
rect 40771 30051 40829 30052
rect 0 29948 80 30028
rect 40003 29968 40012 30008
rect 40052 29968 40780 30008
rect 40820 29968 42796 30008
rect 42836 29968 42845 30008
rect 59308 29924 59348 30052
rect 61228 30008 61268 30220
rect 63532 30176 63572 30220
rect 71299 30176 71357 30177
rect 71692 30176 71732 30220
rect 72451 30219 72509 30220
rect 76099 30219 76157 30220
rect 77251 30219 77309 30220
rect 63340 30136 63572 30176
rect 70915 30136 70924 30176
rect 70964 30136 71308 30176
rect 71348 30136 71732 30176
rect 72067 30136 72076 30176
rect 72116 30136 72268 30176
rect 72308 30136 72317 30176
rect 63340 30092 63380 30136
rect 71299 30135 71357 30136
rect 63235 30052 63244 30092
rect 63284 30052 63380 30092
rect 69475 30052 69484 30092
rect 69524 30052 70540 30092
rect 70580 30052 70589 30092
rect 70723 30052 70732 30092
rect 70772 30052 75436 30092
rect 75476 30052 75485 30092
rect 75811 30052 75820 30092
rect 75860 30052 75869 30092
rect 71107 30008 71165 30009
rect 59395 29968 59404 30008
rect 59444 29968 63340 30008
rect 63380 29968 63389 30008
rect 69283 29968 69292 30008
rect 69332 29968 71116 30008
rect 71156 29968 73460 30008
rect 71107 29967 71165 29968
rect 73420 29924 73460 29968
rect 75820 29924 75860 30052
rect 48931 29884 48940 29924
rect 48980 29884 49516 29924
rect 49556 29884 49940 29924
rect 54787 29884 54796 29924
rect 54836 29884 55180 29924
rect 55220 29884 57004 29924
rect 57044 29884 57053 29924
rect 59308 29884 61420 29924
rect 61460 29884 63380 29924
rect 41443 29800 41452 29840
rect 41492 29800 42316 29840
rect 42356 29800 42365 29840
rect 44515 29800 44524 29840
rect 44564 29800 44812 29840
rect 44852 29800 47788 29840
rect 47828 29800 47837 29840
rect 49219 29800 49228 29840
rect 49268 29800 49708 29840
rect 49748 29800 49757 29840
rect 49900 29756 49940 29884
rect 63340 29840 63380 29884
rect 70540 29884 71980 29924
rect 72020 29884 72029 29924
rect 73420 29884 75052 29924
rect 75092 29884 75101 29924
rect 75619 29884 75628 29924
rect 75668 29884 75860 29924
rect 70540 29840 70580 29884
rect 49987 29800 49996 29840
rect 50036 29800 50476 29840
rect 50516 29800 50668 29840
rect 50708 29800 50717 29840
rect 52483 29800 52492 29840
rect 52532 29800 54124 29840
rect 54164 29800 54173 29840
rect 54979 29800 54988 29840
rect 55028 29800 56428 29840
rect 56468 29800 56716 29840
rect 56756 29800 56765 29840
rect 58819 29800 58828 29840
rect 58868 29800 59788 29840
rect 59828 29800 59837 29840
rect 63340 29800 63436 29840
rect 63476 29800 63485 29840
rect 63907 29800 63916 29840
rect 63956 29800 64780 29840
rect 64820 29800 64829 29840
rect 65443 29800 65452 29840
rect 65492 29800 65836 29840
rect 65876 29800 68332 29840
rect 68372 29800 68381 29840
rect 69091 29800 69100 29840
rect 69140 29800 70540 29840
rect 70580 29800 70589 29840
rect 71011 29800 71020 29840
rect 71060 29800 71404 29840
rect 71444 29800 71453 29840
rect 71779 29800 71788 29840
rect 71828 29800 72076 29840
rect 72116 29800 72125 29840
rect 75523 29800 75532 29840
rect 75572 29800 76012 29840
rect 76052 29800 76061 29840
rect 71299 29756 71357 29757
rect 75820 29756 75860 29800
rect 41347 29716 41356 29756
rect 41396 29716 42124 29756
rect 42164 29716 42173 29756
rect 49891 29716 49900 29756
rect 49940 29716 49949 29756
rect 59491 29716 59500 29756
rect 59540 29716 60172 29756
rect 60212 29716 60221 29756
rect 68227 29716 68236 29756
rect 68276 29716 70924 29756
rect 70964 29716 70973 29756
rect 71214 29716 71308 29756
rect 71348 29716 71357 29756
rect 75811 29716 75820 29756
rect 75860 29716 75900 29756
rect 71299 29715 71357 29716
rect 50563 29632 50572 29672
rect 50612 29632 51532 29672
rect 51572 29632 53644 29672
rect 53684 29632 54316 29672
rect 54356 29632 54365 29672
rect 60067 29632 60076 29672
rect 60116 29632 61324 29672
rect 61364 29632 63052 29672
rect 63092 29632 63101 29672
rect 67651 29632 67660 29672
rect 67700 29632 69964 29672
rect 70004 29632 70013 29672
rect 74851 29632 74860 29672
rect 74900 29632 75916 29672
rect 75956 29632 77260 29672
rect 77300 29632 77309 29672
rect 45667 29548 45676 29588
rect 45716 29548 53300 29588
rect 54979 29548 54988 29588
rect 55028 29548 55468 29588
rect 55508 29548 55660 29588
rect 55700 29548 55709 29588
rect 59203 29548 59212 29588
rect 59252 29548 60268 29588
rect 60308 29548 63532 29588
rect 63572 29548 63581 29588
rect 69763 29548 69772 29588
rect 69812 29548 70252 29588
rect 70292 29548 70301 29588
rect 53260 29504 53300 29548
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 16343 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 16729 29504
rect 28343 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 28729 29504
rect 40343 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 40729 29504
rect 52343 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 52729 29504
rect 53260 29464 57580 29504
rect 57620 29464 57629 29504
rect 60451 29464 60460 29504
rect 60500 29464 60844 29504
rect 60884 29464 60893 29504
rect 61603 29464 61612 29504
rect 61652 29464 64204 29504
rect 64244 29464 64253 29504
rect 64343 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 64729 29504
rect 70051 29464 70060 29504
rect 70100 29464 70636 29504
rect 70676 29464 70685 29504
rect 76343 29464 76352 29504
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76720 29464 76729 29504
rect 46051 29380 46060 29420
rect 46100 29380 46348 29420
rect 46388 29380 48940 29420
rect 48980 29380 57196 29420
rect 57236 29380 57245 29420
rect 70915 29380 70924 29420
rect 70964 29380 72268 29420
rect 72308 29380 72556 29420
rect 72596 29380 72605 29420
rect 55075 29296 55084 29336
rect 55124 29296 55276 29336
rect 55316 29296 55756 29336
rect 55796 29296 55805 29336
rect 63427 29296 63436 29336
rect 63476 29296 64012 29336
rect 64052 29296 64061 29336
rect 65635 29296 65644 29336
rect 65684 29296 66796 29336
rect 66836 29296 66845 29336
rect 71875 29296 71884 29336
rect 71924 29296 76684 29336
rect 76724 29296 77068 29336
rect 77108 29296 77117 29336
rect 61027 29212 61036 29252
rect 61076 29212 61708 29252
rect 61748 29212 61757 29252
rect 63043 29212 63052 29252
rect 63092 29212 68428 29252
rect 68468 29212 68477 29252
rect 75811 29212 75820 29252
rect 75860 29212 76492 29252
rect 76532 29212 76541 29252
rect 0 29108 80 29188
rect 64003 29168 64061 29169
rect 40867 29128 40876 29168
rect 40916 29128 41356 29168
rect 41396 29128 41405 29168
rect 41635 29128 41644 29168
rect 41684 29128 42028 29168
rect 42068 29128 42077 29168
rect 42307 29128 42316 29168
rect 42356 29128 42892 29168
rect 42932 29128 43852 29168
rect 43892 29128 43901 29168
rect 54115 29128 54124 29168
rect 54164 29128 57388 29168
rect 57428 29128 57437 29168
rect 60643 29128 60652 29168
rect 60692 29128 61228 29168
rect 61268 29128 61277 29168
rect 63918 29128 64012 29168
rect 64052 29128 64204 29168
rect 64244 29128 64253 29168
rect 64771 29128 64780 29168
rect 64820 29128 65836 29168
rect 65876 29128 65885 29168
rect 70435 29128 70444 29168
rect 70484 29128 70732 29168
rect 70772 29128 70781 29168
rect 71491 29128 71500 29168
rect 71540 29128 72460 29168
rect 72500 29128 72509 29168
rect 64003 29127 64061 29128
rect 42115 29044 42124 29084
rect 42164 29044 42173 29084
rect 52291 29044 52300 29084
rect 52340 29044 53260 29084
rect 53300 29044 53309 29084
rect 60547 29044 60556 29084
rect 60596 29044 60940 29084
rect 60980 29044 60989 29084
rect 70051 29044 70060 29084
rect 70100 29044 70540 29084
rect 70580 29044 70589 29084
rect 71107 29044 71116 29084
rect 71156 29044 71980 29084
rect 72020 29044 73228 29084
rect 73268 29044 73277 29084
rect 40195 28960 40204 29000
rect 40244 28960 41740 29000
rect 41780 28960 41789 29000
rect 41347 28876 41356 28916
rect 41396 28876 41548 28916
rect 41588 28876 41597 28916
rect 42124 28832 42164 29044
rect 43555 28960 43564 29000
rect 43604 28960 45100 29000
rect 45140 28960 45149 29000
rect 49795 28960 49804 29000
rect 49844 28960 50380 29000
rect 50420 28960 50429 29000
rect 67459 28960 67468 29000
rect 67508 28960 68044 29000
rect 68084 28960 68093 29000
rect 70243 28960 70252 29000
rect 70292 28960 71308 29000
rect 71348 28960 76108 29000
rect 76148 28960 76157 29000
rect 70819 28876 70828 28916
rect 70868 28876 71212 28916
rect 71252 28876 71884 28916
rect 71924 28876 71933 28916
rect 71395 28832 71453 28833
rect 41251 28792 41260 28832
rect 41300 28792 42164 28832
rect 42508 28792 43468 28832
rect 43508 28792 50956 28832
rect 50996 28792 51005 28832
rect 54691 28792 54700 28832
rect 54740 28792 55468 28832
rect 55508 28792 55517 28832
rect 65059 28792 65068 28832
rect 65108 28792 65548 28832
rect 65588 28792 66316 28832
rect 66356 28792 66365 28832
rect 68323 28792 68332 28832
rect 68372 28792 71404 28832
rect 71444 28792 71453 28832
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 15103 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 15489 28748
rect 27103 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 27489 28748
rect 39103 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 39489 28748
rect 40099 28708 40108 28748
rect 40148 28708 42412 28748
rect 42452 28708 42461 28748
rect 42508 28664 42548 28792
rect 71395 28791 71453 28792
rect 77827 28748 77885 28749
rect 49987 28708 49996 28748
rect 50036 28708 50420 28748
rect 51103 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 51489 28748
rect 54883 28708 54892 28748
rect 54932 28708 55564 28748
rect 55604 28708 55613 28748
rect 55939 28708 55948 28748
rect 55988 28708 56428 28748
rect 56468 28708 56477 28748
rect 63103 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 63489 28748
rect 75103 28708 75112 28748
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75480 28708 75489 28748
rect 77742 28708 77836 28748
rect 77876 28708 77885 28748
rect 41731 28624 41740 28664
rect 41780 28624 42548 28664
rect 50380 28580 50420 28708
rect 77827 28707 77885 28708
rect 51340 28624 55276 28664
rect 55316 28624 55325 28664
rect 56899 28624 56908 28664
rect 56948 28624 58540 28664
rect 58580 28624 66892 28664
rect 66932 28624 66941 28664
rect 76771 28624 76780 28664
rect 76820 28624 77068 28664
rect 77108 28624 77117 28664
rect 50467 28580 50525 28581
rect 51340 28580 51380 28624
rect 54595 28580 54653 28581
rect 59395 28580 59453 28581
rect 38467 28540 38476 28580
rect 38516 28540 41068 28580
rect 41108 28540 41117 28580
rect 41443 28540 41452 28580
rect 41492 28540 41836 28580
rect 41876 28540 41885 28580
rect 44611 28540 44620 28580
rect 44660 28540 45388 28580
rect 45428 28540 45437 28580
rect 50380 28540 50476 28580
rect 50516 28540 51340 28580
rect 51380 28540 51389 28580
rect 54510 28540 54604 28580
rect 54644 28540 59404 28580
rect 59444 28540 59453 28580
rect 60835 28540 60844 28580
rect 60884 28540 61516 28580
rect 61556 28540 61565 28580
rect 73411 28540 73420 28580
rect 73460 28540 75340 28580
rect 75380 28540 75389 28580
rect 50467 28539 50525 28540
rect 54595 28539 54653 28540
rect 59395 28539 59453 28540
rect 64003 28496 64061 28497
rect 65155 28496 65213 28497
rect 41923 28456 41932 28496
rect 41972 28456 42316 28496
rect 42356 28456 42365 28496
rect 50179 28456 50188 28496
rect 50228 28456 51724 28496
rect 51764 28456 51773 28496
rect 52867 28456 52876 28496
rect 52916 28456 54508 28496
rect 54548 28456 54557 28496
rect 59299 28456 59308 28496
rect 59348 28456 64012 28496
rect 64052 28456 64061 28496
rect 65070 28456 65164 28496
rect 65204 28456 65213 28496
rect 64003 28455 64061 28456
rect 65155 28455 65213 28456
rect 45763 28372 45772 28412
rect 45812 28372 45821 28412
rect 61219 28372 61228 28412
rect 61268 28372 61612 28412
rect 61652 28372 61661 28412
rect 70540 28372 71692 28412
rect 71732 28372 73804 28412
rect 73844 28372 73853 28412
rect 76387 28372 76396 28412
rect 76436 28372 77492 28412
rect 0 28268 80 28348
rect 39715 28288 39724 28328
rect 39764 28288 40492 28328
rect 40532 28288 41396 28328
rect 43555 28288 43564 28328
rect 43604 28288 44908 28328
rect 44948 28288 45100 28328
rect 45140 28288 45149 28328
rect 41356 28160 41396 28288
rect 45100 28160 45140 28288
rect 45772 28244 45812 28372
rect 46627 28328 46685 28329
rect 60163 28328 60221 28329
rect 70540 28328 70580 28372
rect 77452 28328 77492 28372
rect 45859 28288 45868 28328
rect 45908 28288 46444 28328
rect 46484 28288 46493 28328
rect 46627 28288 46636 28328
rect 46676 28288 46770 28328
rect 49987 28288 49996 28328
rect 50036 28288 50476 28328
rect 50516 28288 50525 28328
rect 50755 28288 50764 28328
rect 50804 28288 51244 28328
rect 51284 28288 51293 28328
rect 55651 28288 55660 28328
rect 55700 28288 56908 28328
rect 56948 28288 56957 28328
rect 59107 28288 59116 28328
rect 59156 28288 59692 28328
rect 59732 28288 59741 28328
rect 60078 28288 60172 28328
rect 60212 28288 60221 28328
rect 60355 28288 60364 28328
rect 60404 28288 60748 28328
rect 60788 28288 60797 28328
rect 61795 28288 61804 28328
rect 61844 28288 63148 28328
rect 63188 28288 63380 28328
rect 64771 28288 64780 28328
rect 64820 28288 64829 28328
rect 66787 28288 66796 28328
rect 66836 28288 66988 28328
rect 67028 28288 67372 28328
rect 67412 28288 67421 28328
rect 70531 28288 70540 28328
rect 70580 28288 70589 28328
rect 75427 28288 75436 28328
rect 75476 28288 76876 28328
rect 76916 28288 76925 28328
rect 77443 28288 77452 28328
rect 77492 28288 78124 28328
rect 78164 28288 79468 28328
rect 79508 28288 79517 28328
rect 46627 28287 46685 28288
rect 60163 28287 60221 28288
rect 45772 28204 46732 28244
rect 46772 28204 47308 28244
rect 47348 28204 47357 28244
rect 50563 28204 50572 28244
rect 50612 28204 50956 28244
rect 50996 28204 54892 28244
rect 54932 28204 54941 28244
rect 50659 28160 50717 28161
rect 63340 28160 63380 28288
rect 64780 28244 64820 28288
rect 63811 28204 63820 28244
rect 63860 28204 64300 28244
rect 64340 28204 64820 28244
rect 41347 28120 41356 28160
rect 41396 28120 41405 28160
rect 45100 28120 46636 28160
rect 46676 28120 46685 28160
rect 48835 28120 48844 28160
rect 48884 28120 50092 28160
rect 50132 28120 50141 28160
rect 50574 28120 50668 28160
rect 50708 28120 50717 28160
rect 52003 28120 52012 28160
rect 52052 28120 53164 28160
rect 53204 28120 53213 28160
rect 55363 28120 55372 28160
rect 55412 28120 56044 28160
rect 56084 28120 56093 28160
rect 57955 28120 57964 28160
rect 58004 28120 58732 28160
rect 58772 28120 59884 28160
rect 59924 28120 59933 28160
rect 63340 28120 65260 28160
rect 65300 28120 65309 28160
rect 70627 28120 70636 28160
rect 70676 28120 70828 28160
rect 70868 28120 70877 28160
rect 50659 28119 50717 28120
rect 52099 28076 52157 28077
rect 71683 28076 71741 28077
rect 44803 28036 44812 28076
rect 44852 28036 46060 28076
rect 46100 28036 47596 28076
rect 47636 28036 47645 28076
rect 52099 28036 52108 28076
rect 52148 28036 58924 28076
rect 58964 28036 59788 28076
rect 59828 28036 59837 28076
rect 60451 28036 60460 28076
rect 60500 28036 60844 28076
rect 60884 28036 60893 28076
rect 65059 28036 65068 28076
rect 65108 28036 65740 28076
rect 65780 28036 65789 28076
rect 68131 28036 68140 28076
rect 68180 28036 71692 28076
rect 71732 28036 71741 28076
rect 45676 27992 45716 28036
rect 46732 27992 46772 28036
rect 52099 28035 52157 28036
rect 71683 28035 71741 28036
rect 52771 27992 52829 27993
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 16343 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 16729 27992
rect 28343 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 28729 27992
rect 40343 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 40729 27992
rect 44707 27952 44716 27992
rect 44756 27952 45484 27992
rect 45524 27952 45533 27992
rect 45667 27952 45676 27992
rect 45716 27952 45756 27992
rect 46723 27952 46732 27992
rect 46772 27952 46812 27992
rect 51523 27952 51532 27992
rect 51572 27952 52012 27992
rect 52052 27952 52061 27992
rect 52343 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 52729 27992
rect 52771 27952 52780 27992
rect 52820 27952 61420 27992
rect 61460 27952 61469 27992
rect 64343 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 64729 27992
rect 65155 27952 65164 27992
rect 65204 27952 65644 27992
rect 65684 27952 65693 27992
rect 65923 27952 65932 27992
rect 65972 27952 66124 27992
rect 66164 27952 66173 27992
rect 76343 27952 76352 27992
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76720 27952 76729 27992
rect 52771 27951 52829 27952
rect 44611 27868 44620 27908
rect 44660 27868 53300 27908
rect 55459 27868 55468 27908
rect 55508 27868 55852 27908
rect 55892 27868 55901 27908
rect 60067 27868 60076 27908
rect 60116 27868 60364 27908
rect 60404 27868 60413 27908
rect 68899 27868 68908 27908
rect 68948 27868 69484 27908
rect 69524 27868 69533 27908
rect 70531 27868 70540 27908
rect 70580 27868 71500 27908
rect 71540 27868 71549 27908
rect 53260 27824 53300 27868
rect 41539 27784 41548 27824
rect 41588 27784 44332 27824
rect 44372 27784 53204 27824
rect 53260 27784 59596 27824
rect 59636 27784 59645 27824
rect 59875 27784 59884 27824
rect 59924 27784 60116 27824
rect 61891 27784 61900 27824
rect 61940 27784 63916 27824
rect 63956 27784 63965 27824
rect 64867 27784 64876 27824
rect 64916 27784 65876 27824
rect 69379 27784 69388 27824
rect 69428 27784 69437 27824
rect 53164 27740 53204 27784
rect 37795 27700 37804 27740
rect 37844 27700 40492 27740
rect 40532 27700 40541 27740
rect 47395 27700 47404 27740
rect 47444 27700 47692 27740
rect 47732 27700 47741 27740
rect 51619 27700 51628 27740
rect 51668 27700 52012 27740
rect 52052 27700 52061 27740
rect 53164 27700 57236 27740
rect 57283 27700 57292 27740
rect 57332 27700 59980 27740
rect 60020 27700 60029 27740
rect 57196 27656 57236 27700
rect 58243 27656 58301 27657
rect 60076 27656 60116 27784
rect 65836 27656 65876 27784
rect 43171 27616 43180 27656
rect 43220 27616 44716 27656
rect 44756 27616 45100 27656
rect 45140 27616 47980 27656
rect 48020 27616 48652 27656
rect 48692 27616 50092 27656
rect 50132 27616 53293 27656
rect 53333 27616 53342 27656
rect 54787 27616 54796 27656
rect 54836 27616 56428 27656
rect 56468 27616 56477 27656
rect 57196 27616 58252 27656
rect 58292 27616 58301 27656
rect 58243 27615 58301 27616
rect 59980 27616 60116 27656
rect 63811 27616 63820 27656
rect 63860 27616 64876 27656
rect 64916 27616 65356 27656
rect 65396 27616 65405 27656
rect 65827 27616 65836 27656
rect 65876 27616 68140 27656
rect 68180 27616 68189 27656
rect 41059 27572 41117 27573
rect 46339 27572 46397 27573
rect 40195 27532 40204 27572
rect 40244 27532 40253 27572
rect 40974 27532 41068 27572
rect 41108 27532 46348 27572
rect 46388 27532 46397 27572
rect 46531 27532 46540 27572
rect 46580 27532 47788 27572
rect 47828 27532 49516 27572
rect 49556 27532 49565 27572
rect 50563 27532 50572 27572
rect 50612 27532 55180 27572
rect 55220 27532 56812 27572
rect 56852 27532 56861 27572
rect 0 27428 80 27508
rect 40204 27320 40244 27532
rect 41059 27531 41117 27532
rect 46339 27531 46397 27532
rect 52003 27488 52061 27489
rect 52771 27488 52829 27489
rect 42787 27448 42796 27488
rect 42836 27448 52012 27488
rect 52052 27448 52780 27488
rect 52820 27448 52829 27488
rect 53284 27448 53293 27488
rect 53333 27448 55372 27488
rect 55412 27448 55421 27488
rect 57100 27448 59924 27488
rect 52003 27447 52061 27448
rect 52771 27447 52829 27448
rect 43075 27404 43133 27405
rect 41635 27364 41644 27404
rect 41684 27364 43084 27404
rect 43124 27364 43133 27404
rect 43075 27363 43133 27364
rect 50755 27404 50813 27405
rect 57100 27404 57140 27448
rect 50755 27364 50764 27404
rect 50804 27364 57140 27404
rect 50755 27363 50813 27364
rect 39715 27280 39724 27320
rect 39764 27280 44524 27320
rect 44564 27280 44908 27320
rect 44948 27280 44957 27320
rect 54883 27280 54892 27320
rect 54932 27280 55181 27320
rect 55221 27280 55230 27320
rect 58051 27280 58060 27320
rect 58100 27280 58828 27320
rect 58868 27280 58877 27320
rect 59884 27236 59924 27448
rect 59980 27320 60020 27616
rect 67555 27572 67613 27573
rect 65443 27532 65452 27572
rect 65492 27532 65740 27572
rect 65780 27532 65789 27572
rect 67470 27532 67564 27572
rect 67604 27532 67613 27572
rect 67555 27531 67613 27532
rect 69388 27488 69428 27784
rect 69484 27740 69524 27868
rect 70060 27784 71924 27824
rect 70060 27740 70100 27784
rect 69484 27700 70060 27740
rect 70100 27700 70109 27740
rect 70243 27700 70252 27740
rect 70292 27700 71500 27740
rect 71540 27700 71549 27740
rect 69763 27616 69772 27656
rect 69812 27616 71788 27656
rect 71828 27616 71837 27656
rect 60163 27448 60172 27488
rect 60212 27448 60652 27488
rect 60692 27448 60701 27488
rect 68323 27448 68332 27488
rect 68372 27448 68908 27488
rect 68948 27448 68957 27488
rect 69388 27448 69772 27488
rect 69812 27448 69821 27488
rect 60163 27404 60221 27405
rect 60067 27364 60076 27404
rect 60116 27364 60172 27404
rect 60212 27364 60221 27404
rect 65251 27364 65260 27404
rect 65300 27364 66796 27404
rect 66836 27364 66845 27404
rect 68515 27364 68524 27404
rect 68564 27364 70252 27404
rect 70292 27364 70301 27404
rect 60163 27363 60221 27364
rect 65155 27320 65213 27321
rect 70828 27320 70868 27616
rect 71884 27404 71924 27784
rect 75235 27700 75244 27740
rect 75284 27700 75436 27740
rect 75476 27700 75485 27740
rect 73507 27616 73516 27656
rect 73556 27616 73900 27656
rect 73940 27616 73949 27656
rect 75043 27616 75052 27656
rect 75092 27616 76780 27656
rect 76820 27616 76972 27656
rect 77012 27616 77021 27656
rect 71971 27488 72029 27489
rect 71971 27448 71980 27488
rect 72020 27448 77164 27488
rect 77204 27448 77213 27488
rect 71971 27447 72029 27448
rect 71299 27364 71308 27404
rect 71348 27364 71596 27404
rect 71636 27364 71645 27404
rect 71884 27364 74092 27404
rect 74132 27364 75244 27404
rect 75284 27364 75293 27404
rect 71395 27320 71453 27321
rect 59980 27280 65012 27320
rect 65070 27280 65164 27320
rect 65204 27280 65213 27320
rect 70819 27280 70828 27320
rect 70868 27280 70877 27320
rect 71310 27280 71404 27320
rect 71444 27280 71453 27320
rect 64972 27236 65012 27280
rect 65155 27279 65213 27280
rect 71395 27279 71453 27280
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 15103 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 15489 27236
rect 27103 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 27489 27236
rect 39103 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 39489 27236
rect 40579 27196 40588 27236
rect 40628 27196 41068 27236
rect 41108 27196 41117 27236
rect 51103 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 51489 27236
rect 51811 27196 51820 27236
rect 51860 27196 52108 27236
rect 52148 27196 52157 27236
rect 59884 27196 60460 27236
rect 60500 27196 61132 27236
rect 61172 27196 61181 27236
rect 63103 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 63489 27236
rect 64972 27196 68812 27236
rect 68852 27196 69004 27236
rect 69044 27196 69053 27236
rect 40195 27152 40253 27153
rect 52963 27152 53021 27153
rect 39148 27112 40204 27152
rect 40244 27112 44620 27152
rect 44660 27112 44669 27152
rect 52963 27112 52972 27152
rect 53012 27112 59020 27152
rect 59060 27112 59069 27152
rect 60739 27112 60748 27152
rect 60788 27112 61036 27152
rect 61076 27112 61085 27152
rect 39148 27068 39188 27112
rect 40195 27111 40253 27112
rect 52963 27111 53021 27112
rect 58531 27068 58589 27069
rect 74956 27068 74996 27364
rect 75103 27196 75112 27236
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75480 27196 75489 27236
rect 39139 27028 39148 27068
rect 39188 27028 39197 27068
rect 39907 27028 39916 27068
rect 39956 27028 40204 27068
rect 40244 27028 40876 27068
rect 40916 27028 40925 27068
rect 54211 27028 54220 27068
rect 54260 27028 55468 27068
rect 55508 27028 55660 27068
rect 55700 27028 55709 27068
rect 58446 27028 58540 27068
rect 58580 27028 58589 27068
rect 58531 27027 58589 27028
rect 58828 27028 61900 27068
rect 61940 27028 61949 27068
rect 74956 27028 75148 27068
rect 75188 27028 75197 27068
rect 75331 27028 75340 27068
rect 75380 27028 75628 27068
rect 75668 27028 75677 27068
rect 50467 26984 50525 26985
rect 50659 26984 50717 26985
rect 58828 26984 58868 27028
rect 50389 26944 50398 26984
rect 50438 26944 50476 26984
rect 50516 26944 50533 26984
rect 50659 26944 50668 26984
rect 50708 26944 55756 26984
rect 55796 26944 55805 26984
rect 58147 26944 58156 26984
rect 58196 26944 58828 26984
rect 58868 26944 58877 26984
rect 59203 26944 59212 26984
rect 59252 26944 63628 26984
rect 63668 26944 64204 26984
rect 64244 26944 64253 26984
rect 75715 26944 75724 26984
rect 75764 26944 75804 26984
rect 50467 26943 50525 26944
rect 50659 26943 50717 26944
rect 40771 26900 40829 26901
rect 58339 26900 58397 26901
rect 60355 26900 60413 26901
rect 75724 26900 75764 26944
rect 39331 26860 39340 26900
rect 39380 26860 39532 26900
rect 39572 26860 40780 26900
rect 40820 26860 40829 26900
rect 40963 26860 40972 26900
rect 41012 26860 41452 26900
rect 41492 26860 41501 26900
rect 58254 26860 58348 26900
rect 58388 26860 58397 26900
rect 60270 26860 60364 26900
rect 60404 26860 60413 26900
rect 60739 26860 60748 26900
rect 60788 26860 64012 26900
rect 64052 26860 64061 26900
rect 73027 26860 73036 26900
rect 73076 26860 74860 26900
rect 74900 26860 74909 26900
rect 75427 26860 75436 26900
rect 75476 26860 75956 26900
rect 40771 26859 40829 26860
rect 58339 26859 58397 26860
rect 60355 26859 60413 26860
rect 40003 26816 40061 26817
rect 60748 26816 60788 26860
rect 75916 26816 75956 26860
rect 39918 26776 40012 26816
rect 40052 26776 40061 26816
rect 43075 26776 43084 26816
rect 43124 26776 43564 26816
rect 43604 26776 43613 26816
rect 46819 26776 46828 26816
rect 46868 26776 47308 26816
rect 47348 26776 52972 26816
rect 53012 26776 53021 26816
rect 55939 26776 55948 26816
rect 55988 26776 56332 26816
rect 56372 26776 56381 26816
rect 57667 26776 57676 26816
rect 57716 26776 59020 26816
rect 59060 26776 59069 26816
rect 60259 26776 60268 26816
rect 60308 26776 60788 26816
rect 61891 26776 61900 26816
rect 61940 26776 62860 26816
rect 62900 26776 63820 26816
rect 63860 26776 63869 26816
rect 66403 26776 66412 26816
rect 66452 26776 67660 26816
rect 67700 26776 67709 26816
rect 68419 26776 68428 26816
rect 68468 26776 68908 26816
rect 68948 26776 68957 26816
rect 74755 26776 74764 26816
rect 74804 26776 75628 26816
rect 75668 26776 75677 26816
rect 75907 26776 75916 26816
rect 75956 26776 76588 26816
rect 76628 26776 76637 26816
rect 40003 26775 40061 26776
rect 41155 26732 41213 26733
rect 39043 26692 39052 26732
rect 39092 26692 41164 26732
rect 41204 26692 41213 26732
rect 41155 26691 41213 26692
rect 53164 26692 54412 26732
rect 54452 26692 54700 26732
rect 54740 26692 54749 26732
rect 55468 26692 58060 26732
rect 58100 26692 58109 26732
rect 60547 26692 60556 26732
rect 60596 26692 72364 26732
rect 72404 26692 72413 26732
rect 0 26588 80 26668
rect 53164 26648 53204 26692
rect 55468 26648 55508 26692
rect 40483 26608 40492 26648
rect 40532 26608 40541 26648
rect 40771 26608 40780 26648
rect 40820 26608 41548 26648
rect 41588 26608 44140 26648
rect 44180 26608 44189 26648
rect 50275 26608 50284 26648
rect 50324 26608 50764 26648
rect 50804 26608 50813 26648
rect 51427 26608 51436 26648
rect 51476 26608 52204 26648
rect 52244 26608 53204 26648
rect 53260 26608 55508 26648
rect 55555 26608 55564 26648
rect 55604 26608 58540 26648
rect 58580 26608 58828 26648
rect 58868 26608 58877 26648
rect 58924 26608 61324 26648
rect 61364 26608 61373 26648
rect 61603 26608 61612 26648
rect 61652 26608 70444 26648
rect 70484 26608 70493 26648
rect 70915 26608 70924 26648
rect 70964 26608 71980 26648
rect 72020 26608 76204 26648
rect 76244 26608 76253 26648
rect 76483 26608 76492 26648
rect 76532 26608 77356 26648
rect 77396 26608 78508 26648
rect 78548 26608 79468 26648
rect 79508 26608 79517 26648
rect 40492 26564 40532 26608
rect 50764 26564 50804 26608
rect 53059 26564 53117 26565
rect 53260 26564 53300 26608
rect 58924 26564 58964 26608
rect 71971 26564 72029 26565
rect 75628 26564 75668 26608
rect 40492 26524 40820 26564
rect 50764 26524 52012 26564
rect 52052 26524 52061 26564
rect 53059 26524 53068 26564
rect 53108 26524 53300 26564
rect 54412 26524 58964 26564
rect 59779 26524 59788 26564
rect 59828 26524 60940 26564
rect 60980 26524 62956 26564
rect 62996 26524 63380 26564
rect 64003 26524 64012 26564
rect 64052 26524 65548 26564
rect 65588 26524 65932 26564
rect 65972 26524 65981 26564
rect 67747 26524 67756 26564
rect 67796 26524 68044 26564
rect 68084 26524 68093 26564
rect 68803 26524 68812 26564
rect 68852 26524 71980 26564
rect 72020 26524 72029 26564
rect 75619 26524 75628 26564
rect 75668 26524 75708 26564
rect 40780 26480 40820 26524
rect 53059 26523 53117 26524
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 16343 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 16729 26480
rect 28343 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 28729 26480
rect 40343 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 40729 26480
rect 40771 26440 40780 26480
rect 40820 26440 40829 26480
rect 52343 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 52729 26480
rect 54412 26396 54452 26524
rect 54499 26480 54557 26481
rect 54499 26440 54508 26480
rect 54548 26440 60556 26480
rect 60596 26440 60605 26480
rect 61123 26440 61132 26480
rect 61172 26440 61612 26480
rect 61652 26440 61661 26480
rect 54499 26439 54557 26440
rect 63340 26396 63380 26524
rect 71971 26523 72029 26524
rect 64343 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 64729 26480
rect 67267 26440 67276 26480
rect 67316 26440 69388 26480
rect 69428 26440 72556 26480
rect 72596 26440 72605 26480
rect 76343 26440 76352 26480
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76720 26440 76729 26480
rect 34915 26356 34924 26396
rect 34964 26356 35404 26396
rect 35444 26356 38092 26396
rect 38132 26356 46060 26396
rect 46100 26356 46109 26396
rect 49507 26356 49516 26396
rect 49556 26356 54452 26396
rect 54604 26356 56044 26396
rect 56084 26356 56093 26396
rect 63340 26356 68428 26396
rect 68468 26356 68477 26396
rect 69484 26356 74764 26396
rect 74804 26356 75724 26396
rect 75764 26356 75773 26396
rect 38947 26312 39005 26313
rect 54604 26312 54644 26356
rect 64003 26312 64061 26313
rect 38947 26272 38956 26312
rect 38996 26272 39052 26312
rect 39092 26272 39101 26312
rect 40579 26272 40588 26312
rect 40628 26272 42028 26312
rect 42068 26272 42077 26312
rect 51139 26272 51148 26312
rect 51188 26272 52108 26312
rect 52148 26272 54644 26312
rect 54691 26272 54700 26312
rect 54740 26272 63532 26312
rect 63572 26272 63581 26312
rect 64003 26272 64012 26312
rect 64052 26272 64396 26312
rect 64436 26272 64445 26312
rect 67843 26272 67852 26312
rect 67892 26272 69004 26312
rect 69044 26272 69053 26312
rect 38947 26271 39005 26272
rect 64003 26271 64061 26272
rect 69484 26228 69524 26356
rect 71299 26272 71308 26312
rect 71348 26272 71596 26312
rect 71636 26272 71645 26312
rect 71779 26272 71788 26312
rect 71828 26272 71837 26312
rect 74467 26272 74476 26312
rect 74516 26272 74668 26312
rect 74708 26272 74717 26312
rect 76867 26272 76876 26312
rect 76916 26272 77068 26312
rect 77108 26272 77117 26312
rect 33475 26188 33484 26228
rect 33524 26188 34252 26228
rect 34292 26188 35020 26228
rect 35060 26188 35069 26228
rect 41644 26188 47020 26228
rect 47060 26188 47069 26228
rect 48835 26188 48844 26228
rect 48884 26188 51532 26228
rect 51572 26188 51581 26228
rect 52003 26188 52012 26228
rect 52052 26188 52492 26228
rect 52532 26188 57676 26228
rect 57716 26188 57725 26228
rect 60355 26188 60364 26228
rect 60404 26188 61132 26228
rect 61172 26188 61181 26228
rect 61603 26188 61612 26228
rect 61652 26188 64780 26228
rect 64820 26188 64829 26228
rect 67363 26188 67372 26228
rect 67412 26188 69484 26228
rect 69524 26188 69533 26228
rect 41644 26144 41684 26188
rect 52195 26144 52253 26145
rect 59395 26144 59453 26145
rect 32707 26104 32716 26144
rect 32756 26104 33964 26144
rect 34004 26104 34013 26144
rect 34339 26104 34348 26144
rect 34388 26104 34732 26144
rect 34772 26104 34781 26144
rect 39427 26104 39436 26144
rect 39476 26104 40300 26144
rect 40340 26104 40349 26144
rect 41059 26104 41068 26144
rect 41108 26104 41452 26144
rect 41492 26104 41501 26144
rect 41635 26104 41644 26144
rect 41684 26104 41693 26144
rect 45379 26104 45388 26144
rect 45428 26104 45964 26144
rect 46004 26104 47788 26144
rect 47828 26104 48940 26144
rect 48980 26104 49132 26144
rect 49172 26104 49181 26144
rect 50659 26104 50668 26144
rect 50708 26104 51724 26144
rect 51764 26104 51773 26144
rect 52195 26104 52204 26144
rect 52244 26104 55564 26144
rect 55604 26104 55613 26144
rect 58627 26104 58636 26144
rect 58676 26104 58924 26144
rect 58964 26104 58973 26144
rect 59310 26104 59404 26144
rect 59444 26104 59453 26144
rect 52195 26103 52253 26104
rect 59395 26103 59453 26104
rect 60364 26104 60460 26144
rect 60500 26104 60509 26144
rect 61411 26104 61420 26144
rect 61460 26104 61804 26144
rect 61844 26104 62860 26144
rect 62900 26104 62909 26144
rect 63811 26104 63820 26144
rect 63860 26104 65356 26144
rect 65396 26104 65405 26144
rect 65635 26104 65644 26144
rect 65684 26104 67180 26144
rect 67220 26104 67229 26144
rect 68611 26104 68620 26144
rect 68660 26104 69292 26144
rect 69332 26104 71308 26144
rect 71348 26104 71357 26144
rect 60364 26061 60404 26104
rect 38851 26060 38909 26061
rect 40867 26060 40925 26061
rect 60355 26060 60413 26061
rect 60547 26060 60605 26061
rect 71788 26060 71828 26272
rect 72547 26188 72556 26228
rect 72596 26188 74860 26228
rect 74900 26188 75820 26228
rect 75860 26188 75869 26228
rect 71971 26104 71980 26144
rect 72020 26104 73460 26144
rect 74275 26104 74284 26144
rect 74324 26104 75916 26144
rect 75956 26104 76396 26144
rect 76436 26104 76445 26144
rect 7180 26020 38092 26060
rect 38132 26020 38141 26060
rect 38766 26020 38860 26060
rect 38900 26020 38909 26060
rect 40387 26020 40396 26060
rect 40436 26020 40876 26060
rect 40916 26020 40925 26060
rect 44899 26020 44908 26060
rect 44948 26020 46444 26060
rect 46484 26020 46493 26060
rect 54979 26020 54988 26060
rect 55028 26020 55037 26060
rect 59299 26020 59308 26060
rect 59348 26020 59924 26060
rect 7180 25976 7220 26020
rect 38851 26019 38909 26020
rect 40867 26019 40925 26020
rect 46819 25976 46877 25977
rect 54988 25976 55028 26020
rect 835 25936 844 25976
rect 884 25936 7220 25976
rect 31939 25936 31948 25976
rect 31988 25936 33484 25976
rect 33524 25936 33533 25976
rect 34627 25936 34636 25976
rect 34676 25936 36748 25976
rect 36788 25936 36797 25976
rect 39331 25936 39340 25976
rect 39380 25936 40204 25976
rect 40244 25936 40253 25976
rect 46339 25936 46348 25976
rect 46388 25936 46828 25976
rect 46868 25936 46877 25976
rect 47395 25936 47404 25976
rect 47444 25936 49228 25976
rect 49268 25936 49277 25976
rect 50947 25936 50956 25976
rect 50996 25936 51820 25976
rect 51860 25936 55028 25976
rect 55075 25936 55084 25976
rect 55124 25936 55660 25976
rect 55700 25936 56524 25976
rect 56564 25936 56573 25976
rect 57475 25936 57484 25976
rect 57524 25936 58348 25976
rect 58388 25936 58397 25976
rect 58531 25936 58540 25976
rect 58580 25936 59212 25976
rect 59252 25936 59788 25976
rect 59828 25936 59837 25976
rect 46819 25935 46877 25936
rect 59395 25892 59453 25893
rect 33139 25852 33148 25892
rect 33188 25852 33580 25892
rect 33620 25852 33629 25892
rect 37219 25852 37228 25892
rect 37268 25852 39244 25892
rect 39284 25852 39293 25892
rect 40771 25852 40780 25892
rect 40820 25852 41740 25892
rect 41780 25852 41789 25892
rect 44803 25852 44812 25892
rect 44852 25852 46252 25892
rect 46292 25852 46540 25892
rect 46580 25852 46732 25892
rect 46772 25852 46781 25892
rect 51235 25852 51244 25892
rect 51284 25852 51724 25892
rect 51764 25852 51773 25892
rect 52675 25852 52684 25892
rect 52724 25852 54796 25892
rect 54836 25852 54845 25892
rect 58435 25852 58444 25892
rect 58484 25852 59404 25892
rect 59444 25852 59453 25892
rect 59884 25892 59924 26020
rect 60355 26020 60364 26060
rect 60404 26020 60413 26060
rect 60462 26020 60556 26060
rect 60596 26020 60605 26060
rect 60739 26020 60748 26060
rect 60788 26020 71828 26060
rect 73420 26060 73460 26104
rect 73420 26020 75860 26060
rect 60355 26019 60413 26020
rect 60547 26019 60605 26020
rect 75820 25976 75860 26020
rect 64291 25936 64300 25976
rect 64340 25936 64780 25976
rect 64820 25936 64829 25976
rect 64963 25936 64972 25976
rect 65012 25936 65356 25976
rect 65396 25936 65405 25976
rect 73219 25936 73228 25976
rect 73268 25936 74476 25976
rect 74516 25936 74525 25976
rect 74851 25936 74860 25976
rect 74900 25936 75436 25976
rect 75476 25936 75628 25976
rect 75668 25936 75677 25976
rect 75811 25936 75820 25976
rect 75860 25936 76684 25976
rect 76724 25936 76733 25976
rect 77827 25892 77885 25893
rect 59884 25852 60364 25892
rect 60404 25852 61516 25892
rect 61556 25852 61565 25892
rect 67843 25852 67852 25892
rect 67892 25852 68236 25892
rect 68276 25852 68285 25892
rect 72643 25852 72652 25892
rect 72692 25852 74380 25892
rect 74420 25852 74429 25892
rect 76195 25852 76204 25892
rect 76244 25852 76780 25892
rect 76820 25852 76829 25892
rect 77742 25852 77836 25892
rect 77876 25852 77885 25892
rect 59395 25851 59453 25852
rect 77827 25851 77885 25852
rect 0 25808 80 25828
rect 0 25768 652 25808
rect 692 25768 701 25808
rect 35203 25768 35212 25808
rect 35252 25768 35788 25808
rect 35828 25768 35837 25808
rect 46051 25768 46060 25808
rect 46100 25768 57964 25808
rect 58004 25768 58013 25808
rect 58819 25768 58828 25808
rect 58868 25768 60748 25808
rect 60788 25768 60797 25808
rect 0 25748 80 25768
rect 41155 25724 41213 25725
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 15103 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 15489 25724
rect 27103 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 27489 25724
rect 39103 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 39489 25724
rect 41155 25684 41164 25724
rect 41204 25684 49420 25724
rect 49460 25684 49996 25724
rect 50036 25684 50045 25724
rect 51103 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 51489 25724
rect 58147 25684 58156 25724
rect 58196 25684 59020 25724
rect 59060 25684 59069 25724
rect 63103 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 63489 25724
rect 65059 25684 65068 25724
rect 65108 25684 68140 25724
rect 68180 25684 68189 25724
rect 75103 25684 75112 25724
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75480 25684 75489 25724
rect 41155 25683 41213 25684
rect 63907 25640 63965 25641
rect 38083 25600 38092 25640
rect 38132 25600 43220 25640
rect 43843 25600 43852 25640
rect 43892 25600 44044 25640
rect 44084 25600 44093 25640
rect 44140 25600 52876 25640
rect 52916 25600 52925 25640
rect 60163 25600 60172 25640
rect 60212 25600 63916 25640
rect 63956 25600 63965 25640
rect 41059 25556 41117 25557
rect 35011 25516 35020 25556
rect 35060 25516 35692 25556
rect 35732 25516 35741 25556
rect 40483 25516 40492 25556
rect 40532 25516 40876 25556
rect 40916 25516 41068 25556
rect 41108 25516 41117 25556
rect 43180 25556 43220 25600
rect 44140 25556 44180 25600
rect 63907 25599 63965 25600
rect 43180 25516 44180 25556
rect 44323 25516 44332 25556
rect 44372 25516 59020 25556
rect 59060 25516 59069 25556
rect 41059 25515 41117 25516
rect 44227 25432 44236 25472
rect 44276 25432 46348 25472
rect 46388 25432 46397 25472
rect 50563 25432 50572 25472
rect 50612 25432 51724 25472
rect 51764 25432 51773 25472
rect 71203 25432 71212 25472
rect 71252 25432 71788 25472
rect 71828 25432 72844 25472
rect 72884 25432 73036 25472
rect 73076 25432 73085 25472
rect 35491 25348 35500 25388
rect 35540 25348 35884 25388
rect 35924 25348 35933 25388
rect 40675 25348 40684 25388
rect 40724 25348 43220 25388
rect 44611 25348 44620 25388
rect 44660 25348 45292 25388
rect 45332 25348 45341 25388
rect 45388 25348 60940 25388
rect 60980 25348 60989 25388
rect 63340 25348 66316 25388
rect 66356 25348 67084 25388
rect 67124 25348 67133 25388
rect 75427 25348 75436 25388
rect 75476 25348 75724 25388
rect 75764 25348 75773 25388
rect 33187 25264 33196 25304
rect 33236 25264 35692 25304
rect 35732 25264 35741 25304
rect 36355 25264 36364 25304
rect 36404 25264 36940 25304
rect 36980 25264 38476 25304
rect 38516 25264 38956 25304
rect 38996 25264 39005 25304
rect 34636 25136 34676 25264
rect 39907 25180 39916 25220
rect 39956 25180 39965 25220
rect 39916 25136 39956 25180
rect 40003 25136 40061 25137
rect 43180 25136 43220 25348
rect 44323 25264 44332 25304
rect 44372 25264 45004 25304
rect 45044 25264 45053 25304
rect 45388 25220 45428 25348
rect 46147 25304 46205 25305
rect 46627 25304 46685 25305
rect 50659 25304 50717 25305
rect 63340 25304 63380 25348
rect 46147 25264 46156 25304
rect 46196 25264 46444 25304
rect 46484 25264 46636 25304
rect 46676 25264 46685 25304
rect 50179 25264 50188 25304
rect 50228 25264 50668 25304
rect 50708 25264 50717 25304
rect 51811 25264 51820 25304
rect 51860 25264 52684 25304
rect 52724 25264 52733 25304
rect 55459 25264 55468 25304
rect 55508 25264 55756 25304
rect 55796 25264 57004 25304
rect 57044 25264 57053 25304
rect 59587 25264 59596 25304
rect 59636 25264 63148 25304
rect 63188 25264 63380 25304
rect 63427 25264 63436 25304
rect 63476 25264 63916 25304
rect 63956 25264 63965 25304
rect 66787 25264 66796 25304
rect 66836 25264 69196 25304
rect 69236 25264 70348 25304
rect 70388 25264 71884 25304
rect 71924 25264 72652 25304
rect 72692 25264 72701 25304
rect 74467 25264 74476 25304
rect 74516 25264 77932 25304
rect 77972 25264 78316 25304
rect 78356 25264 78365 25304
rect 46147 25263 46205 25264
rect 46627 25263 46685 25264
rect 50659 25263 50717 25264
rect 51619 25220 51677 25221
rect 45283 25180 45292 25220
rect 45332 25180 45428 25220
rect 46636 25180 51628 25220
rect 51668 25180 51677 25220
rect 52003 25180 52012 25220
rect 52052 25180 52396 25220
rect 52436 25180 52445 25220
rect 53260 25180 74572 25220
rect 74612 25180 74621 25220
rect 76291 25180 76300 25220
rect 76340 25180 76684 25220
rect 76724 25180 76733 25220
rect 46636 25136 46676 25180
rect 51340 25136 51380 25180
rect 51619 25179 51677 25180
rect 53260 25136 53300 25180
rect 60355 25136 60413 25137
rect 835 25096 844 25136
rect 884 25096 2764 25136
rect 2804 25096 2813 25136
rect 34627 25096 34636 25136
rect 34676 25096 34685 25136
rect 35875 25096 35884 25136
rect 35924 25096 36460 25136
rect 36500 25096 36844 25136
rect 36884 25096 36893 25136
rect 39916 25096 40012 25136
rect 40052 25096 40108 25136
rect 40148 25096 40157 25136
rect 43180 25096 46676 25136
rect 46723 25096 46732 25136
rect 46772 25096 49556 25136
rect 51331 25096 51340 25136
rect 51380 25096 51389 25136
rect 51907 25096 51916 25136
rect 51956 25096 53300 25136
rect 58051 25096 58060 25136
rect 58100 25096 58828 25136
rect 58868 25096 58877 25136
rect 59395 25096 59404 25136
rect 59444 25096 59884 25136
rect 59924 25096 59933 25136
rect 60355 25096 60364 25136
rect 60404 25096 60460 25136
rect 60500 25096 60509 25136
rect 61507 25096 61516 25136
rect 61556 25096 63532 25136
rect 63572 25096 65068 25136
rect 65108 25096 65117 25136
rect 70339 25096 70348 25136
rect 70388 25096 72460 25136
rect 72500 25096 72509 25136
rect 40003 25095 40061 25096
rect 49516 25052 49556 25096
rect 60355 25095 60413 25096
rect 63907 25052 63965 25053
rect 46819 25012 46828 25052
rect 46868 25012 47500 25052
rect 47540 25012 47549 25052
rect 49507 25012 49516 25052
rect 49556 25012 61708 25052
rect 61748 25012 61757 25052
rect 63907 25012 63916 25052
rect 63956 25012 66700 25052
rect 66740 25012 66749 25052
rect 67651 25012 67660 25052
rect 67700 25012 67852 25052
rect 67892 25012 67901 25052
rect 63907 25011 63965 25012
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 16343 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 16729 24968
rect 28343 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 28729 24968
rect 40343 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 40729 24968
rect 51811 24928 51820 24968
rect 51860 24928 52108 24968
rect 52148 24928 52157 24968
rect 52343 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 52729 24968
rect 54787 24928 54796 24968
rect 54836 24928 63436 24968
rect 63476 24928 63485 24968
rect 64343 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 64729 24968
rect 66403 24928 66412 24968
rect 66452 24928 72076 24968
rect 72116 24928 72125 24968
rect 73420 24928 76204 24968
rect 76244 24928 76253 24968
rect 76343 24928 76352 24968
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76720 24928 76729 24968
rect 0 24908 80 24928
rect 73420 24884 73460 24928
rect 47107 24844 47116 24884
rect 47156 24844 47165 24884
rect 50947 24844 50956 24884
rect 50996 24844 58636 24884
rect 58676 24844 58685 24884
rect 58915 24844 58924 24884
rect 58964 24844 59596 24884
rect 59636 24844 59645 24884
rect 59779 24844 59788 24884
rect 59828 24844 60172 24884
rect 60212 24844 60221 24884
rect 63907 24844 63916 24884
rect 63956 24844 64148 24884
rect 70531 24844 70540 24884
rect 70580 24844 73460 24884
rect 35971 24760 35980 24800
rect 36020 24760 36652 24800
rect 36692 24760 37516 24800
rect 37556 24760 37565 24800
rect 40300 24760 40492 24800
rect 40532 24760 40876 24800
rect 40916 24760 40925 24800
rect 40300 24716 40340 24760
rect 29827 24676 29836 24716
rect 29876 24676 32524 24716
rect 32564 24676 32573 24716
rect 37699 24676 37708 24716
rect 37748 24676 40340 24716
rect 46819 24632 46877 24633
rect 32707 24592 32716 24632
rect 32756 24592 33292 24632
rect 33332 24592 33341 24632
rect 35203 24592 35212 24632
rect 35252 24592 40396 24632
rect 40436 24592 40445 24632
rect 40675 24592 40684 24632
rect 40724 24592 40972 24632
rect 41012 24592 41021 24632
rect 42307 24592 42316 24632
rect 42356 24592 44428 24632
rect 44468 24592 44477 24632
rect 45100 24592 46828 24632
rect 46868 24592 46877 24632
rect 47116 24632 47156 24844
rect 47299 24800 47357 24801
rect 47299 24760 47308 24800
rect 47348 24760 47442 24800
rect 58060 24760 59444 24800
rect 59491 24760 59500 24800
rect 59540 24760 60076 24800
rect 60116 24760 62572 24800
rect 62612 24760 62621 24800
rect 47299 24759 47357 24760
rect 58060 24716 58100 24760
rect 59404 24716 59444 24760
rect 63907 24716 63965 24717
rect 64108 24716 64148 24844
rect 67363 24760 67372 24800
rect 67412 24760 68332 24800
rect 68372 24760 70348 24800
rect 70388 24760 70397 24800
rect 71587 24760 71596 24800
rect 71636 24760 74476 24800
rect 74516 24760 74956 24800
rect 74996 24760 76492 24800
rect 76532 24760 76541 24800
rect 49507 24676 49516 24716
rect 49556 24676 50476 24716
rect 50516 24676 50525 24716
rect 57091 24676 57100 24716
rect 57140 24676 58060 24716
rect 58100 24676 58109 24716
rect 58723 24676 58732 24716
rect 58772 24676 58781 24716
rect 59395 24676 59404 24716
rect 59444 24676 59453 24716
rect 63907 24676 63916 24716
rect 63956 24676 64050 24716
rect 64108 24676 64588 24716
rect 64628 24676 66412 24716
rect 66452 24676 66461 24716
rect 66691 24676 66700 24716
rect 66740 24676 67660 24716
rect 67700 24676 67709 24716
rect 58732 24632 58772 24676
rect 63907 24675 63965 24676
rect 47116 24592 47212 24632
rect 47252 24592 47261 24632
rect 51139 24592 51148 24632
rect 51188 24592 51628 24632
rect 51668 24592 52300 24632
rect 52340 24592 52349 24632
rect 53635 24592 53644 24632
rect 53684 24592 56332 24632
rect 56372 24592 58772 24632
rect 63619 24592 63628 24632
rect 63668 24592 64108 24632
rect 64148 24592 64157 24632
rect 64387 24592 64396 24632
rect 64436 24592 65548 24632
rect 65588 24592 67412 24632
rect 68131 24592 68140 24632
rect 68180 24592 68189 24632
rect 71011 24592 71020 24632
rect 71060 24592 71692 24632
rect 71732 24592 71741 24632
rect 75715 24592 75724 24632
rect 75764 24592 76684 24632
rect 76724 24592 78988 24632
rect 79028 24592 79037 24632
rect 38947 24548 39005 24549
rect 31075 24508 31084 24548
rect 31124 24508 33580 24548
rect 33620 24508 34348 24548
rect 34388 24508 34397 24548
rect 38947 24508 38956 24548
rect 38996 24508 39052 24548
rect 39092 24508 39101 24548
rect 39811 24508 39820 24548
rect 39860 24508 41068 24548
rect 41108 24508 43276 24548
rect 43316 24508 43325 24548
rect 38947 24507 39005 24508
rect 39715 24464 39773 24465
rect 45100 24464 45140 24592
rect 46819 24591 46877 24592
rect 67372 24548 67412 24592
rect 68140 24548 68180 24592
rect 46339 24508 46348 24548
rect 46388 24508 47308 24548
rect 47348 24508 47357 24548
rect 54307 24508 54316 24548
rect 54356 24508 55412 24548
rect 55939 24508 55948 24548
rect 55988 24508 57484 24548
rect 57524 24508 67276 24548
rect 67316 24508 67325 24548
rect 67372 24508 68180 24548
rect 55372 24464 55412 24508
rect 36739 24424 36748 24464
rect 36788 24424 39532 24464
rect 39572 24424 39724 24464
rect 39764 24424 39773 24464
rect 40867 24424 40876 24464
rect 40916 24424 41356 24464
rect 41396 24424 41405 24464
rect 43747 24424 43756 24464
rect 43796 24424 44908 24464
rect 44948 24424 44957 24464
rect 45091 24424 45100 24464
rect 45140 24424 45149 24464
rect 52195 24424 52204 24464
rect 52244 24424 53164 24464
rect 53204 24424 55276 24464
rect 55316 24424 55325 24464
rect 55372 24424 64492 24464
rect 64532 24424 64541 24464
rect 39715 24423 39773 24424
rect 33187 24340 33196 24380
rect 33236 24340 33388 24380
rect 33428 24340 34580 24380
rect 39235 24340 39244 24380
rect 39284 24340 40108 24380
rect 40148 24340 40157 24380
rect 44227 24340 44236 24380
rect 44276 24340 44716 24380
rect 44756 24340 45196 24380
rect 45236 24340 45484 24380
rect 45524 24340 45533 24380
rect 49795 24340 49804 24380
rect 49844 24340 50188 24380
rect 50228 24340 50237 24380
rect 50371 24340 50380 24380
rect 50420 24340 50860 24380
rect 50900 24340 50909 24380
rect 34540 24296 34580 24340
rect 47299 24296 47357 24297
rect 31747 24256 31756 24296
rect 31796 24256 32332 24296
rect 32372 24256 34444 24296
rect 34484 24256 34493 24296
rect 34540 24256 39628 24296
rect 39668 24256 39677 24296
rect 41155 24256 41164 24296
rect 41204 24256 43852 24296
rect 43892 24256 43901 24296
rect 47107 24256 47116 24296
rect 47156 24256 47308 24296
rect 47348 24256 47357 24296
rect 48547 24256 48556 24296
rect 48596 24256 62476 24296
rect 62516 24256 62525 24296
rect 47299 24255 47357 24256
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 15103 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 15489 24212
rect 27103 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 27489 24212
rect 39103 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 39489 24212
rect 44035 24172 44044 24212
rect 44084 24172 44332 24212
rect 44372 24172 44524 24212
rect 44564 24172 44573 24212
rect 46243 24172 46252 24212
rect 46292 24172 46924 24212
rect 46964 24172 46973 24212
rect 73123 24172 73132 24212
rect 73172 24172 75244 24212
rect 75284 24172 75293 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 35491 24088 35500 24128
rect 35540 24088 57676 24128
rect 57716 24088 57725 24128
rect 0 24068 80 24088
rect 1795 24004 1804 24044
rect 1844 24004 2188 24044
rect 2228 24004 35060 24044
rect 35107 24004 35116 24044
rect 35156 24004 35884 24044
rect 35924 24004 35933 24044
rect 45379 24004 45388 24044
rect 45428 24004 48844 24044
rect 48884 24004 62092 24044
rect 62132 24004 62141 24044
rect 62563 24004 62572 24044
rect 62612 24004 67756 24044
rect 67796 24004 67805 24044
rect 73891 24004 73900 24044
rect 73940 24004 74476 24044
rect 74516 24004 74525 24044
rect 35020 23960 35060 24004
rect 51331 23960 51389 23961
rect 31843 23920 31852 23960
rect 31892 23920 32812 23960
rect 32852 23920 34540 23960
rect 34580 23920 34589 23960
rect 35020 23920 41164 23960
rect 41204 23920 41213 23960
rect 44131 23920 44140 23960
rect 44180 23920 44620 23960
rect 44660 23920 44669 23960
rect 47683 23920 47692 23960
rect 47732 23920 48364 23960
rect 48404 23920 49228 23960
rect 49268 23920 49277 23960
rect 49891 23920 49900 23960
rect 49940 23920 50764 23960
rect 50804 23920 50813 23960
rect 51043 23920 51052 23960
rect 51092 23920 51340 23960
rect 51380 23920 51389 23960
rect 52195 23920 52204 23960
rect 52244 23920 52253 23960
rect 57187 23920 57196 23960
rect 57236 23920 60844 23960
rect 60884 23920 61228 23960
rect 61268 23920 61277 23960
rect 63235 23920 63244 23960
rect 63284 23920 63293 23960
rect 65251 23920 65260 23960
rect 65300 23920 65644 23960
rect 65684 23920 66028 23960
rect 66068 23920 66077 23960
rect 68515 23920 68524 23960
rect 68564 23920 68908 23960
rect 68948 23920 68957 23960
rect 70147 23920 70156 23960
rect 70196 23920 70540 23960
rect 70580 23920 70828 23960
rect 70868 23920 70877 23960
rect 73315 23920 73324 23960
rect 73364 23920 73612 23960
rect 73652 23920 73804 23960
rect 73844 23920 73853 23960
rect 73987 23920 73996 23960
rect 74036 23920 74860 23960
rect 74900 23920 74909 23960
rect 51331 23919 51389 23920
rect 52204 23876 52244 23920
rect 835 23836 844 23876
rect 884 23836 1996 23876
rect 2036 23836 2045 23876
rect 29539 23836 29548 23876
rect 29588 23836 31468 23876
rect 31508 23836 36556 23876
rect 36596 23836 36605 23876
rect 51052 23836 52244 23876
rect 57571 23836 57580 23876
rect 57620 23836 60460 23876
rect 60500 23836 60748 23876
rect 60788 23836 60797 23876
rect 51052 23792 51092 23836
rect 54787 23792 54845 23793
rect 55843 23792 55901 23793
rect 56803 23792 56861 23793
rect 57283 23792 57341 23793
rect 63244 23792 63284 23920
rect 70627 23792 70685 23793
rect 71683 23792 71741 23793
rect 76099 23792 76157 23793
rect 76963 23792 77021 23793
rect 77443 23792 77501 23793
rect 79075 23792 79133 23793
rect 32323 23752 32332 23792
rect 32372 23752 33140 23792
rect 34339 23752 34348 23792
rect 34388 23752 36364 23792
rect 36404 23752 36413 23792
rect 37315 23752 37324 23792
rect 37364 23752 43220 23792
rect 43939 23752 43948 23792
rect 43988 23752 44428 23792
rect 44468 23752 44477 23792
rect 44611 23752 44620 23792
rect 44660 23752 46060 23792
rect 46100 23752 46109 23792
rect 49987 23752 49996 23792
rect 50036 23752 50572 23792
rect 50612 23752 50621 23792
rect 51043 23752 51052 23792
rect 51092 23752 51101 23792
rect 52963 23752 52972 23792
rect 53012 23752 53644 23792
rect 53684 23752 53693 23792
rect 54702 23752 54796 23792
rect 54836 23752 54845 23792
rect 55758 23752 55852 23792
rect 55892 23752 56044 23792
rect 56084 23752 56093 23792
rect 56718 23752 56812 23792
rect 56852 23752 56861 23792
rect 57198 23752 57292 23792
rect 57332 23752 57341 23792
rect 59011 23752 59020 23792
rect 59060 23752 59692 23792
rect 59732 23752 59980 23792
rect 60020 23752 60029 23792
rect 63244 23752 64108 23792
rect 64148 23752 64157 23792
rect 67267 23752 67276 23792
rect 67316 23752 67660 23792
rect 67700 23752 67709 23792
rect 68707 23752 68716 23792
rect 68756 23752 70156 23792
rect 70196 23752 70444 23792
rect 70484 23752 70493 23792
rect 70627 23752 70636 23792
rect 70676 23752 70924 23792
rect 70964 23752 70973 23792
rect 71598 23752 71692 23792
rect 71732 23752 71980 23792
rect 72020 23752 72029 23792
rect 76014 23752 76108 23792
rect 76148 23752 76492 23792
rect 76532 23752 76541 23792
rect 76878 23752 76972 23792
rect 77012 23752 77021 23792
rect 77358 23752 77452 23792
rect 77492 23752 77501 23792
rect 78990 23752 79084 23792
rect 79124 23752 79133 23792
rect 33100 23708 33140 23752
rect 43180 23708 43220 23752
rect 54787 23751 54845 23752
rect 55843 23751 55901 23752
rect 56803 23751 56861 23752
rect 57283 23751 57341 23752
rect 70627 23751 70685 23752
rect 71683 23751 71741 23752
rect 76099 23751 76157 23752
rect 76963 23751 77021 23752
rect 77443 23751 77501 23752
rect 79075 23751 79133 23752
rect 51715 23708 51773 23709
rect 31459 23668 31468 23708
rect 31508 23668 32140 23708
rect 32180 23668 32428 23708
rect 32468 23668 32477 23708
rect 33100 23668 33388 23708
rect 33428 23668 35500 23708
rect 35540 23668 35549 23708
rect 38083 23668 38092 23708
rect 38132 23668 38860 23708
rect 38900 23668 38909 23708
rect 40387 23668 40396 23708
rect 40436 23668 40876 23708
rect 40916 23668 40925 23708
rect 43180 23668 51724 23708
rect 51764 23668 51773 23708
rect 51715 23667 51773 23668
rect 51820 23668 54124 23708
rect 54164 23668 63244 23708
rect 63284 23668 63628 23708
rect 63668 23668 63677 23708
rect 46147 23624 46205 23625
rect 51820 23624 51860 23668
rect 58243 23624 58301 23625
rect 60547 23624 60605 23625
rect 835 23584 844 23624
rect 884 23584 1420 23624
rect 1460 23584 1469 23624
rect 33100 23584 34828 23624
rect 34868 23584 37228 23624
rect 37268 23584 37277 23624
rect 46062 23584 46156 23624
rect 46196 23584 46205 23624
rect 47971 23584 47980 23624
rect 48020 23584 50668 23624
rect 50708 23584 50717 23624
rect 50760 23584 50769 23624
rect 50809 23584 51244 23624
rect 51284 23584 51293 23624
rect 51715 23584 51724 23624
rect 51764 23584 51860 23624
rect 53260 23584 57620 23624
rect 57667 23584 57676 23624
rect 57716 23584 58060 23624
rect 58100 23584 58109 23624
rect 58243 23584 58252 23624
rect 58292 23584 60076 23624
rect 60116 23584 60556 23624
rect 60596 23584 60605 23624
rect 62467 23584 62476 23624
rect 62516 23584 62860 23624
rect 62900 23584 62909 23624
rect 68899 23584 68908 23624
rect 68948 23584 69292 23624
rect 69332 23584 69341 23624
rect 75235 23584 75244 23624
rect 75284 23584 75628 23624
rect 75668 23584 75677 23624
rect 33100 23540 33140 23584
rect 46147 23583 46205 23584
rect 53260 23540 53300 23584
rect 56131 23540 56189 23541
rect 32332 23500 33140 23540
rect 34531 23500 34540 23540
rect 34580 23500 35788 23540
rect 35828 23500 39052 23540
rect 39092 23500 39101 23540
rect 43267 23500 43276 23540
rect 43316 23500 53300 23540
rect 56046 23500 56140 23540
rect 56180 23500 56189 23540
rect 57580 23540 57620 23584
rect 58243 23583 58301 23584
rect 60547 23583 60605 23584
rect 57580 23500 59308 23540
rect 59348 23500 59692 23540
rect 59732 23500 59741 23540
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 16343 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 16729 23456
rect 28343 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 28729 23456
rect 32332 23372 32372 23500
rect 56131 23499 56189 23500
rect 54787 23456 54845 23457
rect 56803 23456 56861 23457
rect 34435 23416 34444 23456
rect 34484 23416 36076 23456
rect 36116 23416 38956 23456
rect 38996 23416 39005 23456
rect 40343 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 40729 23456
rect 41731 23416 41740 23456
rect 41780 23416 45100 23456
rect 45140 23416 45149 23456
rect 50563 23416 50572 23456
rect 50612 23416 51724 23456
rect 51764 23416 51773 23456
rect 52396 23416 52876 23456
rect 52916 23416 52925 23456
rect 54787 23416 54796 23456
rect 54836 23416 55276 23456
rect 55316 23416 55325 23456
rect 56803 23416 56812 23456
rect 56852 23416 57292 23456
rect 57332 23416 57341 23456
rect 74851 23416 74860 23456
rect 74900 23416 75244 23456
rect 75284 23416 75293 23456
rect 78787 23416 78796 23456
rect 78836 23416 79276 23456
rect 79316 23416 79325 23456
rect 32323 23332 32332 23372
rect 32372 23332 32381 23372
rect 36163 23332 36172 23372
rect 36212 23332 37900 23372
rect 37940 23332 37949 23372
rect 41251 23332 41260 23372
rect 41300 23332 44812 23372
rect 44852 23332 45004 23372
rect 45044 23332 46540 23372
rect 46580 23332 46589 23372
rect 50371 23332 50380 23372
rect 50420 23332 51820 23372
rect 51860 23332 51869 23372
rect 0 23288 80 23308
rect 52396 23288 52436 23416
rect 54787 23415 54845 23416
rect 56803 23415 56861 23416
rect 52963 23332 52972 23372
rect 53012 23332 62764 23372
rect 62804 23332 63244 23372
rect 63284 23332 63293 23372
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 30979 23248 30988 23288
rect 31028 23248 31276 23288
rect 31316 23248 31325 23288
rect 31939 23248 31948 23288
rect 31988 23248 32716 23288
rect 32756 23248 35212 23288
rect 35252 23248 35261 23288
rect 36931 23248 36940 23288
rect 36980 23248 37132 23288
rect 37172 23248 37181 23288
rect 38851 23248 38860 23288
rect 38900 23248 40876 23288
rect 40916 23248 41356 23288
rect 41396 23248 41405 23288
rect 41827 23248 41836 23288
rect 41876 23248 43756 23288
rect 43796 23248 44620 23288
rect 44660 23248 44669 23288
rect 48643 23248 48652 23288
rect 48692 23248 49804 23288
rect 49844 23248 49853 23288
rect 50755 23248 50764 23288
rect 50804 23248 51052 23288
rect 51092 23248 51101 23288
rect 51427 23248 51436 23288
rect 51476 23248 52436 23288
rect 52483 23288 52541 23289
rect 56803 23288 56861 23289
rect 52483 23248 52492 23288
rect 52532 23248 52588 23288
rect 52628 23248 52637 23288
rect 52684 23248 56372 23288
rect 56419 23248 56428 23288
rect 56468 23248 56812 23288
rect 56852 23248 56861 23288
rect 74467 23248 74476 23288
rect 74516 23248 74860 23288
rect 74900 23248 74909 23288
rect 0 23228 80 23248
rect 44620 23204 44660 23248
rect 52483 23247 52541 23248
rect 52684 23204 52724 23248
rect 55651 23204 55709 23205
rect 1507 23164 1516 23204
rect 1556 23164 2132 23204
rect 28195 23164 28204 23204
rect 28244 23164 30796 23204
rect 30836 23164 30845 23204
rect 31363 23164 31372 23204
rect 31412 23164 31660 23204
rect 31700 23164 32620 23204
rect 32660 23164 33196 23204
rect 33236 23164 33245 23204
rect 36355 23164 36364 23204
rect 36404 23164 37228 23204
rect 37268 23164 37277 23204
rect 37795 23164 37804 23204
rect 37844 23164 38284 23204
rect 38324 23164 39340 23204
rect 39380 23164 39389 23204
rect 44620 23164 46732 23204
rect 46772 23164 46781 23204
rect 48739 23164 48748 23204
rect 48788 23164 49900 23204
rect 49940 23164 49949 23204
rect 50467 23164 50476 23204
rect 50516 23164 50668 23204
rect 50708 23164 50717 23204
rect 51811 23164 51820 23204
rect 51860 23164 52724 23204
rect 52867 23164 52876 23204
rect 52916 23164 54316 23204
rect 54356 23164 54365 23204
rect 55075 23164 55084 23204
rect 55124 23164 55660 23204
rect 55700 23164 55709 23204
rect 56332 23204 56372 23248
rect 56803 23247 56861 23248
rect 56332 23164 58444 23204
rect 58484 23164 58828 23204
rect 58868 23164 58877 23204
rect 2092 23120 2132 23164
rect 46051 23120 46109 23121
rect 50476 23120 50516 23164
rect 55651 23163 55709 23164
rect 51331 23120 51389 23121
rect 1411 23080 1420 23120
rect 1460 23080 1900 23120
rect 1940 23080 1949 23120
rect 2083 23080 2092 23120
rect 2132 23080 3628 23120
rect 3668 23080 3820 23120
rect 3860 23080 3869 23120
rect 32419 23080 32428 23120
rect 32468 23080 32812 23120
rect 32852 23080 32861 23120
rect 32995 23080 33004 23120
rect 33044 23080 33292 23120
rect 33332 23080 33341 23120
rect 35875 23080 35884 23120
rect 35924 23080 36076 23120
rect 36116 23080 36125 23120
rect 36259 23080 36268 23120
rect 36308 23080 36748 23120
rect 36788 23080 36797 23120
rect 37027 23080 37036 23120
rect 37076 23080 39724 23120
rect 39764 23080 40012 23120
rect 40052 23080 42124 23120
rect 42164 23080 42173 23120
rect 45571 23080 45580 23120
rect 45620 23080 45868 23120
rect 45908 23080 45917 23120
rect 46051 23080 46060 23120
rect 46100 23080 46156 23120
rect 46196 23080 46205 23120
rect 49699 23080 49708 23120
rect 49748 23080 50516 23120
rect 51246 23080 51340 23120
rect 51380 23080 51389 23120
rect 52675 23080 52684 23120
rect 52724 23080 54785 23120
rect 46051 23079 46109 23080
rect 51331 23079 51389 23080
rect 54745 23036 54785 23080
rect 56131 23036 56189 23037
rect 22051 22996 22060 23036
rect 22100 22996 42412 23036
rect 42452 22996 45292 23036
rect 45332 22996 45341 23036
rect 50179 22996 50188 23036
rect 50228 22996 51532 23036
rect 51572 22996 51581 23036
rect 52291 22996 52300 23036
rect 52340 22996 54055 23036
rect 54095 22996 54104 23036
rect 54736 22996 54745 23036
rect 54785 22996 54825 23036
rect 56131 22996 56140 23036
rect 56180 22996 56455 23036
rect 56495 22996 56504 23036
rect 44140 22952 44180 22996
rect 56131 22995 56189 22996
rect 36451 22912 36460 22952
rect 36500 22912 37996 22952
rect 38036 22912 38045 22952
rect 41443 22912 41452 22952
rect 41492 22912 42028 22952
rect 42068 22912 42077 22952
rect 44131 22912 44140 22952
rect 44180 22912 44220 22952
rect 52771 22912 52780 22952
rect 52820 22912 53545 22952
rect 53585 22912 53594 22952
rect 54691 22868 54749 22869
rect 40195 22828 40204 22868
rect 40244 22828 42604 22868
rect 42644 22828 42988 22868
rect 43028 22828 43037 22868
rect 52003 22828 52012 22868
rect 52052 22828 53655 22868
rect 53695 22828 53704 22868
rect 54691 22828 54700 22868
rect 54740 22828 54855 22868
rect 54895 22828 54904 22868
rect 54691 22827 54749 22828
rect 54403 22784 54461 22785
rect 57667 22784 57725 22785
rect 60547 22784 60605 22785
rect 43171 22744 43180 22784
rect 43220 22744 51820 22784
rect 51860 22744 51869 22784
rect 52387 22744 52396 22784
rect 52436 22744 53945 22784
rect 53985 22744 53994 22784
rect 54360 22744 54412 22784
rect 54452 22744 54455 22784
rect 54495 22744 54504 22784
rect 57581 22744 57655 22784
rect 57716 22744 57725 22784
rect 59011 22744 59020 22784
rect 59060 22744 59255 22784
rect 59295 22744 59304 22784
rect 60455 22744 60464 22784
rect 60504 22744 60556 22784
rect 60596 22744 60605 22784
rect 78595 22744 78604 22784
rect 78644 22744 78855 22784
rect 78895 22744 78904 22784
rect 54403 22743 54461 22744
rect 57667 22743 57725 22744
rect 60547 22743 60605 22744
rect 46147 22700 46205 22701
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 15103 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 15489 22700
rect 27103 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 27489 22700
rect 30787 22660 30796 22700
rect 30836 22660 31852 22700
rect 31892 22660 32716 22700
rect 32756 22660 32765 22700
rect 39103 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 39489 22700
rect 41539 22660 41548 22700
rect 41588 22660 43468 22700
rect 43508 22660 43517 22700
rect 46062 22660 46156 22700
rect 46196 22660 46205 22700
rect 46147 22659 46205 22660
rect 51811 22616 51869 22617
rect 30979 22576 30988 22616
rect 31028 22576 32044 22616
rect 32084 22576 32093 22616
rect 34915 22576 34924 22616
rect 34964 22576 51820 22616
rect 51860 22576 51869 22616
rect 51811 22575 51869 22576
rect 38467 22492 38476 22532
rect 38516 22492 39052 22532
rect 39092 22492 39101 22532
rect 43459 22492 43468 22532
rect 43508 22492 50860 22532
rect 50900 22492 50909 22532
rect 0 22448 80 22468
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 30883 22408 30892 22448
rect 30932 22408 31468 22448
rect 31508 22408 32084 22448
rect 35587 22408 35596 22448
rect 35636 22408 36172 22448
rect 36212 22408 36221 22448
rect 36643 22408 36652 22448
rect 36692 22408 36844 22448
rect 36884 22408 38188 22448
rect 38228 22408 43084 22448
rect 43124 22408 43133 22448
rect 0 22388 80 22408
rect 1891 22324 1900 22364
rect 1940 22324 3244 22364
rect 3284 22324 3293 22364
rect 32044 22280 32084 22408
rect 40387 22324 40396 22364
rect 40436 22324 40588 22364
rect 40628 22324 41644 22364
rect 41684 22324 41693 22364
rect 42979 22324 42988 22364
rect 43028 22324 49036 22364
rect 49076 22324 49085 22364
rect 29635 22240 29644 22280
rect 29684 22240 30316 22280
rect 30356 22240 31276 22280
rect 31316 22240 31325 22280
rect 32035 22240 32044 22280
rect 32084 22240 32093 22280
rect 39235 22240 39244 22280
rect 39284 22240 40780 22280
rect 40820 22240 40829 22280
rect 42115 22240 42124 22280
rect 42164 22240 42316 22280
rect 42356 22240 43564 22280
rect 43604 22240 43613 22280
rect 45379 22240 45388 22280
rect 45428 22240 46252 22280
rect 46292 22240 46301 22280
rect 46627 22240 46636 22280
rect 46676 22240 48556 22280
rect 48596 22240 48605 22280
rect 48931 22240 48940 22280
rect 48980 22240 51436 22280
rect 51476 22240 51485 22280
rect 52099 22240 52108 22280
rect 52148 22240 52684 22280
rect 52724 22240 52733 22280
rect 38851 22196 38909 22197
rect 52291 22196 52349 22197
rect 27523 22156 27532 22196
rect 27572 22156 28012 22196
rect 28052 22156 38860 22196
rect 38900 22156 38909 22196
rect 50275 22156 50284 22196
rect 50324 22156 50860 22196
rect 50900 22156 50909 22196
rect 52206 22156 52300 22196
rect 52340 22156 52349 22196
rect 38851 22155 38909 22156
rect 52291 22155 52349 22156
rect 27907 22072 27916 22112
rect 27956 22072 28204 22112
rect 28244 22072 30412 22112
rect 30452 22072 31756 22112
rect 31796 22072 32908 22112
rect 32948 22072 32957 22112
rect 49219 22072 49228 22112
rect 49268 22072 50764 22112
rect 50804 22072 50813 22112
rect 32035 21988 32044 22028
rect 32084 21988 32524 22028
rect 32564 21988 32573 22028
rect 45283 21988 45292 22028
rect 45332 21988 46060 22028
rect 46100 21988 46109 22028
rect 50371 21988 50380 22028
rect 50420 21988 52972 22028
rect 53012 21988 53021 22028
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 16343 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 16729 21944
rect 28343 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 28729 21944
rect 28771 21904 28780 21944
rect 28820 21904 29452 21944
rect 29492 21904 29501 21944
rect 40343 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 40729 21944
rect 45571 21904 45580 21944
rect 45620 21904 45629 21944
rect 49507 21904 49516 21944
rect 49556 21904 51148 21944
rect 51188 21904 51197 21944
rect 38851 21860 38909 21861
rect 31171 21820 31180 21860
rect 31220 21820 32044 21860
rect 32084 21820 34924 21860
rect 34964 21820 34973 21860
rect 38851 21820 38860 21860
rect 38900 21820 42988 21860
rect 43028 21820 43037 21860
rect 38851 21819 38909 21820
rect 3235 21736 3244 21776
rect 3284 21736 12980 21776
rect 27619 21736 27628 21776
rect 27668 21736 28012 21776
rect 28052 21736 30508 21776
rect 30548 21736 30557 21776
rect 32140 21736 32332 21776
rect 32372 21736 32381 21776
rect 35779 21736 35788 21776
rect 35828 21736 36268 21776
rect 36308 21736 36317 21776
rect 41059 21736 41068 21776
rect 41108 21736 41260 21776
rect 41300 21736 41309 21776
rect 12940 21692 12980 21736
rect 12940 21652 22252 21692
rect 22292 21652 22301 21692
rect 28387 21652 28396 21692
rect 28436 21652 30892 21692
rect 30932 21652 30941 21692
rect 0 21608 80 21628
rect 32140 21608 32180 21736
rect 41260 21652 41548 21692
rect 41588 21652 41597 21692
rect 42307 21652 42316 21692
rect 42356 21652 45196 21692
rect 45236 21652 45245 21692
rect 41260 21608 41300 21652
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 835 21568 844 21608
rect 884 21568 3052 21608
rect 3092 21568 3101 21608
rect 29059 21568 29068 21608
rect 29108 21568 29548 21608
rect 29588 21568 29597 21608
rect 31459 21568 31468 21608
rect 31508 21568 32180 21608
rect 32995 21568 33004 21608
rect 33044 21568 36172 21608
rect 36212 21568 36221 21608
rect 41251 21568 41260 21608
rect 41300 21568 41309 21608
rect 44899 21568 44908 21608
rect 44948 21568 45388 21608
rect 45428 21568 45437 21608
rect 0 21548 80 21568
rect 45580 21524 45620 21904
rect 50755 21736 50764 21776
rect 50804 21736 51148 21776
rect 51188 21736 51197 21776
rect 99920 21692 100000 21726
rect 50371 21652 50380 21692
rect 50420 21652 51052 21692
rect 51092 21652 51101 21692
rect 99888 21652 100000 21692
rect 52579 21608 52637 21609
rect 49027 21568 49036 21608
rect 49076 21568 49612 21608
rect 49652 21568 50956 21608
rect 50996 21568 51005 21608
rect 52494 21568 52588 21608
rect 52628 21568 52637 21608
rect 99920 21586 100000 21652
rect 52579 21567 52637 21568
rect 2860 21484 5932 21524
rect 5972 21484 5981 21524
rect 25891 21484 25900 21524
rect 25940 21484 26860 21524
rect 26900 21484 32372 21524
rect 39235 21484 39244 21524
rect 39284 21484 40108 21524
rect 40148 21484 42412 21524
rect 42452 21484 42461 21524
rect 45283 21484 45292 21524
rect 45332 21484 48364 21524
rect 48404 21484 48413 21524
rect 2860 21440 2900 21484
rect 931 21400 940 21440
rect 980 21400 2900 21440
rect 3139 21400 3148 21440
rect 3188 21400 3572 21440
rect 5539 21400 5548 21440
rect 5588 21400 12980 21440
rect 26467 21400 26476 21440
rect 26516 21400 27820 21440
rect 27860 21400 27869 21440
rect 3532 21356 3572 21400
rect 12940 21356 12980 21400
rect 1699 21316 1708 21356
rect 1748 21316 2668 21356
rect 2708 21316 3244 21356
rect 3284 21316 3293 21356
rect 3523 21316 3532 21356
rect 3572 21316 4780 21356
rect 4820 21316 4829 21356
rect 5731 21316 5740 21356
rect 5780 21316 6124 21356
rect 6164 21316 6173 21356
rect 12940 21316 22348 21356
rect 22388 21316 27436 21356
rect 27476 21316 27485 21356
rect 26851 21232 26860 21272
rect 26900 21232 31372 21272
rect 31412 21232 31421 21272
rect 32332 21188 32372 21484
rect 39139 21400 39148 21440
rect 39188 21400 39916 21440
rect 39956 21400 42316 21440
rect 42356 21400 44332 21440
rect 44372 21400 45004 21440
rect 45044 21400 45053 21440
rect 38563 21316 38572 21356
rect 38612 21316 39052 21356
rect 39092 21316 39101 21356
rect 45667 21316 45676 21356
rect 45716 21316 45964 21356
rect 46004 21316 46013 21356
rect 47683 21316 47692 21356
rect 47732 21316 48844 21356
rect 48884 21316 48893 21356
rect 51619 21272 51677 21273
rect 32419 21232 32428 21272
rect 32468 21232 51628 21272
rect 51668 21232 51677 21272
rect 51619 21231 51677 21232
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 15103 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 15489 21188
rect 27103 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 27489 21188
rect 32332 21148 38516 21188
rect 39103 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 39489 21188
rect 38476 21104 38516 21148
rect 40195 21104 40253 21105
rect 2851 21064 2860 21104
rect 2900 21064 3628 21104
rect 3668 21064 25900 21104
rect 25940 21064 25949 21104
rect 27340 21064 29356 21104
rect 29396 21064 34636 21104
rect 34676 21064 34685 21104
rect 38476 21064 40204 21104
rect 40244 21064 40253 21104
rect 27340 21020 27380 21064
rect 40195 21063 40253 21064
rect 26659 20980 26668 21020
rect 26708 20980 27380 21020
rect 28867 20980 28876 21020
rect 28916 20980 29068 21020
rect 29108 20980 31660 21020
rect 31700 20980 32428 21020
rect 32468 20980 32477 21020
rect 48547 20980 48556 21020
rect 48596 20980 50092 21020
rect 50132 20980 50141 21020
rect 52291 20936 52349 20937
rect 27619 20896 27628 20936
rect 27668 20896 29260 20936
rect 29300 20896 30508 20936
rect 30548 20896 31180 20936
rect 31220 20896 31229 20936
rect 31852 20896 33004 20936
rect 33044 20896 33053 20936
rect 37123 20896 37132 20936
rect 37172 20896 52300 20936
rect 52340 20896 52349 20936
rect 31852 20852 31892 20896
rect 52291 20895 52349 20896
rect 43075 20852 43133 20853
rect 46051 20852 46109 20853
rect 28003 20812 28012 20852
rect 28052 20812 28684 20852
rect 28724 20812 31852 20852
rect 31892 20812 31901 20852
rect 32131 20812 32140 20852
rect 32180 20812 43084 20852
rect 43124 20812 43660 20852
rect 43700 20812 43709 20852
rect 45475 20812 45484 20852
rect 45524 20812 46060 20852
rect 46100 20812 46109 20852
rect 43075 20811 43133 20812
rect 46051 20811 46109 20812
rect 0 20768 80 20788
rect 40195 20768 40253 20769
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 6115 20728 6124 20768
rect 6164 20728 27380 20768
rect 28483 20728 28492 20768
rect 28532 20728 28876 20768
rect 28916 20728 28925 20768
rect 31171 20728 31180 20768
rect 31220 20728 33580 20768
rect 33620 20728 33629 20768
rect 36643 20728 36652 20768
rect 36692 20728 37420 20768
rect 37460 20728 37469 20768
rect 40195 20728 40204 20768
rect 40244 20728 41740 20768
rect 41780 20728 41789 20768
rect 42403 20728 42412 20768
rect 42452 20728 44620 20768
rect 44660 20728 44908 20768
rect 44948 20728 44957 20768
rect 45667 20728 45676 20768
rect 45716 20728 46060 20768
rect 46100 20728 46109 20768
rect 46339 20728 46348 20768
rect 46388 20728 46732 20768
rect 46772 20728 46781 20768
rect 47203 20728 47212 20768
rect 47252 20728 47596 20768
rect 47636 20728 48940 20768
rect 48980 20728 50860 20768
rect 50900 20728 51532 20768
rect 51572 20728 51581 20768
rect 0 20708 80 20728
rect 27340 20600 27380 20728
rect 40195 20727 40253 20728
rect 27907 20644 27916 20684
rect 27956 20644 28396 20684
rect 28436 20644 28445 20684
rect 28771 20644 28780 20684
rect 28820 20644 29260 20684
rect 29300 20644 29309 20684
rect 27340 20560 33140 20600
rect 40963 20560 40972 20600
rect 41012 20560 41164 20600
rect 41204 20560 41213 20600
rect 33100 20516 33140 20560
rect 33100 20476 41644 20516
rect 41684 20476 41693 20516
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 16343 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 16729 20432
rect 28343 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 28729 20432
rect 34627 20392 34636 20432
rect 34676 20392 35212 20432
rect 35252 20392 38188 20432
rect 38228 20392 38237 20432
rect 40343 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 40729 20432
rect 52483 20264 52541 20265
rect 24067 20224 24076 20264
rect 24116 20224 26956 20264
rect 26996 20224 27244 20264
rect 27284 20224 27628 20264
rect 27668 20224 27677 20264
rect 32035 20224 32044 20264
rect 32084 20224 32093 20264
rect 41155 20224 41164 20264
rect 41204 20224 41932 20264
rect 41972 20224 41981 20264
rect 44803 20224 44812 20264
rect 44852 20224 52492 20264
rect 52532 20224 52541 20264
rect 32044 20180 32084 20224
rect 52483 20223 52541 20224
rect 28195 20140 28204 20180
rect 28244 20140 29068 20180
rect 29108 20140 29117 20180
rect 31747 20140 31756 20180
rect 31796 20140 34828 20180
rect 34868 20140 34877 20180
rect 35011 20140 35020 20180
rect 35060 20140 38036 20180
rect 39619 20140 39628 20180
rect 39668 20140 40972 20180
rect 41012 20140 41021 20180
rect 41443 20140 41452 20180
rect 41492 20140 42124 20180
rect 42164 20140 42173 20180
rect 44995 20140 45004 20180
rect 45044 20140 47596 20180
rect 47636 20140 47645 20180
rect 52579 20140 52588 20180
rect 52628 20140 52637 20180
rect 37996 20096 38036 20140
rect 52588 20096 52628 20140
rect 25795 20056 25804 20096
rect 25844 20056 26956 20096
rect 26996 20056 27724 20096
rect 27764 20056 28300 20096
rect 28340 20056 28349 20096
rect 32899 20056 32908 20096
rect 32948 20056 34732 20096
rect 34772 20056 34924 20096
rect 34964 20056 34973 20096
rect 36259 20056 36268 20096
rect 36308 20056 37804 20096
rect 37844 20056 37853 20096
rect 37987 20056 37996 20096
rect 38036 20056 38045 20096
rect 45187 20056 45196 20096
rect 45236 20056 52628 20096
rect 99920 20012 100000 20089
rect 5539 19972 5548 20012
rect 5588 19972 9004 20012
rect 9044 19972 9053 20012
rect 25603 19972 25612 20012
rect 25652 19972 26284 20012
rect 26324 19972 26764 20012
rect 26804 19972 26813 20012
rect 29059 19972 29068 20012
rect 29108 19972 31468 20012
rect 31508 19972 31517 20012
rect 32227 19972 32236 20012
rect 32276 19972 32285 20012
rect 34819 19972 34828 20012
rect 34868 19972 37228 20012
rect 37268 19972 37277 20012
rect 42883 19972 42892 20012
rect 42932 19972 43276 20012
rect 43316 19972 43325 20012
rect 44515 19972 44524 20012
rect 44564 19972 45292 20012
rect 45332 19972 46636 20012
rect 46676 19972 49324 20012
rect 49364 19972 51628 20012
rect 51668 19972 51677 20012
rect 99888 19972 100000 20012
rect 0 19928 80 19948
rect 32236 19928 32276 19972
rect 99920 19949 100000 19972
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 26851 19888 26860 19928
rect 26900 19888 27340 19928
rect 27380 19888 29164 19928
rect 29204 19888 29213 19928
rect 32236 19888 35020 19928
rect 35060 19888 35069 19928
rect 44131 19888 44140 19928
rect 44180 19888 44716 19928
rect 44756 19888 44765 19928
rect 0 19868 80 19888
rect 47683 19844 47741 19845
rect 22531 19804 22540 19844
rect 22580 19804 22828 19844
rect 22868 19804 22877 19844
rect 32227 19804 32236 19844
rect 32276 19804 32716 19844
rect 32756 19804 33196 19844
rect 33236 19804 33245 19844
rect 37603 19804 37612 19844
rect 37652 19804 38380 19844
rect 38420 19804 38668 19844
rect 38708 19804 38717 19844
rect 43267 19804 43276 19844
rect 43316 19804 43852 19844
rect 43892 19804 43901 19844
rect 47299 19804 47308 19844
rect 47348 19804 47500 19844
rect 47540 19804 47549 19844
rect 47683 19804 47692 19844
rect 47732 19804 47826 19844
rect 47683 19803 47741 19804
rect 32803 19720 32812 19760
rect 32852 19720 33100 19760
rect 33140 19720 33149 19760
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 15103 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 15489 19676
rect 27103 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 27489 19676
rect 32899 19636 32908 19676
rect 32948 19636 33236 19676
rect 39103 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 39489 19676
rect 33196 19592 33236 19636
rect 21955 19552 21964 19592
rect 22004 19552 32140 19592
rect 32180 19552 32189 19592
rect 33187 19552 33196 19592
rect 33236 19552 33245 19592
rect 11683 19508 11741 19509
rect 40867 19508 40925 19509
rect 11598 19468 11692 19508
rect 11732 19468 11741 19508
rect 22147 19468 22156 19508
rect 22196 19468 27916 19508
rect 27956 19468 27965 19508
rect 37507 19468 37516 19508
rect 37556 19468 39052 19508
rect 39092 19468 39101 19508
rect 40867 19468 40876 19508
rect 40916 19468 47020 19508
rect 47060 19468 47069 19508
rect 11683 19467 11741 19468
rect 40867 19467 40925 19468
rect 6595 19384 6604 19424
rect 6644 19384 7948 19424
rect 7988 19384 7997 19424
rect 8803 19384 8812 19424
rect 8852 19384 9292 19424
rect 9332 19384 9341 19424
rect 39139 19384 39148 19424
rect 39188 19384 40684 19424
rect 40724 19384 40733 19424
rect 40195 19340 40253 19341
rect 8515 19300 8524 19340
rect 8564 19300 9004 19340
rect 9044 19300 9053 19340
rect 21571 19300 21580 19340
rect 21620 19300 27628 19340
rect 27668 19300 27677 19340
rect 40195 19300 40204 19340
rect 40244 19300 40300 19340
rect 40340 19300 40349 19340
rect 41251 19300 41260 19340
rect 41300 19300 41836 19340
rect 41876 19300 41885 19340
rect 42508 19300 43276 19340
rect 43316 19300 43325 19340
rect 40195 19299 40253 19300
rect 39715 19256 39773 19257
rect 42508 19256 42548 19300
rect 8611 19216 8620 19256
rect 8660 19216 8669 19256
rect 9091 19216 9100 19256
rect 9140 19216 9484 19256
rect 9524 19216 9533 19256
rect 10531 19216 10540 19256
rect 10580 19216 31084 19256
rect 31124 19216 31133 19256
rect 37027 19216 37036 19256
rect 37076 19216 38188 19256
rect 38228 19216 38237 19256
rect 38947 19216 38956 19256
rect 38996 19216 39724 19256
rect 39764 19216 39773 19256
rect 42499 19216 42508 19256
rect 42548 19216 42557 19256
rect 42691 19216 42700 19256
rect 42740 19216 44332 19256
rect 44372 19216 45004 19256
rect 45044 19216 45053 19256
rect 8620 19172 8660 19216
rect 39715 19215 39773 19216
rect 8620 19132 26668 19172
rect 26708 19132 26717 19172
rect 49123 19132 49132 19172
rect 49172 19132 49612 19172
rect 49652 19132 49661 19172
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 21763 19048 21772 19088
rect 21812 19048 22924 19088
rect 22964 19048 22973 19088
rect 31651 19048 31660 19088
rect 31700 19048 31852 19088
rect 31892 19048 31901 19088
rect 37219 19048 37228 19088
rect 37268 19048 38668 19088
rect 38708 19048 38717 19088
rect 41635 19048 41644 19088
rect 41684 19048 42892 19088
rect 42932 19048 42941 19088
rect 0 19028 80 19048
rect 38371 18964 38380 19004
rect 38420 18964 39436 19004
rect 39476 18964 41204 19004
rect 41164 18920 41204 18964
rect 47395 18920 47453 18921
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 8323 18880 8332 18920
rect 8372 18880 8812 18920
rect 8852 18880 8861 18920
rect 16343 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 16729 18920
rect 22531 18880 22540 18920
rect 22580 18880 22828 18920
rect 22868 18880 22877 18920
rect 28343 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 28729 18920
rect 40343 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 40729 18920
rect 41155 18880 41164 18920
rect 41204 18880 42836 18920
rect 43171 18880 43180 18920
rect 43220 18880 44620 18920
rect 44660 18880 44669 18920
rect 47310 18880 47404 18920
rect 47444 18880 48940 18920
rect 48980 18880 48989 18920
rect 33283 18836 33341 18837
rect 42796 18836 42836 18880
rect 47395 18879 47453 18880
rect 8515 18796 8524 18836
rect 8564 18796 8908 18836
rect 8948 18796 8957 18836
rect 33198 18796 33292 18836
rect 33332 18796 33341 18836
rect 42115 18796 42124 18836
rect 42164 18796 42740 18836
rect 42796 18796 50860 18836
rect 50900 18796 50909 18836
rect 33283 18795 33341 18796
rect 22915 18712 22924 18752
rect 22964 18712 26572 18752
rect 26612 18712 27052 18752
rect 27092 18712 27101 18752
rect 33379 18712 33388 18752
rect 33428 18712 33468 18752
rect 41443 18712 41452 18752
rect 41492 18712 42644 18752
rect 33388 18668 33428 18712
rect 42604 18668 42644 18712
rect 9187 18628 9196 18668
rect 9236 18628 22060 18668
rect 22100 18628 22109 18668
rect 23107 18628 23116 18668
rect 23156 18628 25228 18668
rect 25268 18628 25277 18668
rect 25324 18628 29068 18668
rect 29108 18628 29117 18668
rect 29923 18628 29932 18668
rect 29972 18628 30604 18668
rect 30644 18628 31852 18668
rect 31892 18628 31901 18668
rect 32428 18628 34828 18668
rect 34868 18628 35596 18668
rect 35636 18628 35645 18668
rect 35779 18628 35788 18668
rect 35828 18628 36172 18668
rect 36212 18628 36221 18668
rect 36451 18628 36460 18668
rect 36500 18628 36844 18668
rect 36884 18628 36893 18668
rect 38851 18628 38860 18668
rect 38900 18628 40972 18668
rect 41012 18628 41021 18668
rect 42595 18628 42604 18668
rect 42644 18628 42653 18668
rect 8035 18544 8044 18584
rect 8084 18544 8524 18584
rect 8564 18544 8573 18584
rect 9571 18544 9580 18584
rect 9620 18544 11692 18584
rect 11732 18544 11741 18584
rect 22531 18544 22540 18584
rect 22580 18544 23020 18584
rect 23060 18544 23069 18584
rect 25324 18500 25364 18628
rect 25603 18544 25612 18584
rect 25652 18544 25661 18584
rect 26659 18544 26668 18584
rect 26708 18544 26956 18584
rect 26996 18544 28684 18584
rect 28724 18544 28733 18584
rect 28963 18544 28972 18584
rect 29012 18544 32140 18584
rect 32180 18544 32332 18584
rect 32372 18544 32381 18584
rect 22435 18460 22444 18500
rect 22484 18460 22828 18500
rect 22868 18460 22877 18500
rect 23779 18460 23788 18500
rect 23828 18460 23980 18500
rect 24020 18460 25364 18500
rect 25612 18500 25652 18544
rect 28972 18500 29012 18544
rect 32428 18500 32468 18628
rect 33475 18584 33533 18585
rect 32803 18544 32812 18584
rect 32852 18544 33292 18584
rect 33332 18544 33341 18584
rect 33475 18544 33484 18584
rect 33524 18544 33618 18584
rect 33667 18544 33676 18584
rect 33716 18544 34252 18584
rect 34292 18544 35500 18584
rect 35540 18544 37420 18584
rect 37460 18544 37469 18584
rect 33475 18543 33533 18544
rect 38860 18500 38900 18628
rect 25612 18460 29012 18500
rect 31267 18460 31276 18500
rect 31316 18460 32468 18500
rect 32515 18460 32524 18500
rect 32564 18460 35692 18500
rect 35732 18460 38900 18500
rect 33475 18416 33533 18417
rect 42604 18416 42644 18628
rect 42700 18584 42740 18796
rect 49027 18752 49085 18753
rect 42787 18712 42796 18752
rect 42836 18712 43468 18752
rect 43508 18712 43517 18752
rect 45571 18712 45580 18752
rect 45620 18712 46156 18752
rect 46196 18712 46205 18752
rect 48556 18712 48884 18752
rect 48942 18712 49036 18752
rect 49076 18712 49085 18752
rect 49219 18712 49228 18752
rect 49268 18712 49277 18752
rect 48556 18668 48596 18712
rect 43939 18628 43948 18668
rect 43988 18628 45484 18668
rect 45524 18628 45533 18668
rect 46819 18628 46828 18668
rect 46868 18628 48076 18668
rect 48116 18628 48596 18668
rect 48844 18668 48884 18712
rect 49027 18711 49085 18712
rect 49228 18668 49268 18712
rect 48844 18628 49268 18668
rect 46147 18584 46205 18585
rect 51907 18584 51965 18585
rect 42700 18544 43660 18584
rect 43700 18544 44044 18584
rect 44084 18544 44093 18584
rect 44227 18544 44236 18584
rect 44276 18544 44524 18584
rect 44564 18544 44573 18584
rect 46062 18544 46156 18584
rect 46196 18544 46205 18584
rect 47011 18544 47020 18584
rect 47060 18544 47404 18584
rect 47444 18544 47453 18584
rect 47683 18544 47692 18584
rect 47732 18544 48652 18584
rect 48692 18544 48701 18584
rect 48931 18544 48940 18584
rect 48980 18544 49900 18584
rect 49940 18544 49949 18584
rect 51907 18544 51916 18584
rect 51956 18544 52300 18584
rect 52340 18544 52349 18584
rect 46147 18543 46205 18544
rect 51907 18543 51965 18544
rect 43075 18500 43133 18501
rect 47395 18500 47453 18501
rect 51811 18500 51869 18501
rect 42990 18460 43084 18500
rect 43124 18460 43133 18500
rect 43747 18460 43756 18500
rect 43796 18460 45100 18500
rect 45140 18460 45149 18500
rect 46435 18460 46444 18500
rect 46484 18460 46924 18500
rect 46964 18460 46973 18500
rect 47395 18460 47404 18500
rect 47444 18460 47453 18500
rect 47971 18460 47980 18500
rect 48020 18460 48844 18500
rect 48884 18460 48893 18500
rect 49507 18460 49516 18500
rect 49556 18460 51820 18500
rect 51860 18460 52012 18500
rect 52052 18460 52061 18500
rect 43075 18459 43133 18460
rect 4771 18376 4780 18416
rect 4820 18376 24364 18416
rect 24404 18376 26860 18416
rect 26900 18376 26909 18416
rect 27043 18376 27052 18416
rect 27092 18376 29836 18416
rect 29876 18376 29885 18416
rect 30211 18376 30220 18416
rect 30260 18376 33484 18416
rect 33524 18376 33533 18416
rect 42211 18376 42220 18416
rect 42260 18376 42412 18416
rect 42452 18376 42461 18416
rect 42604 18376 43276 18416
rect 43316 18376 44428 18416
rect 44468 18376 44477 18416
rect 22243 18292 22252 18332
rect 22292 18292 22444 18332
rect 22484 18292 29204 18332
rect 29251 18292 29260 18332
rect 29300 18292 30124 18332
rect 30164 18292 31180 18332
rect 31220 18292 31229 18332
rect 0 18248 80 18268
rect 29164 18248 29204 18292
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 21475 18208 21484 18248
rect 21524 18208 21868 18248
rect 21908 18208 28012 18248
rect 28052 18208 28061 18248
rect 29164 18208 32140 18248
rect 32180 18208 32189 18248
rect 0 18188 80 18208
rect 26467 18164 26525 18165
rect 33100 18164 33140 18376
rect 33475 18375 33533 18376
rect 33283 18332 33341 18333
rect 35395 18332 35453 18333
rect 44524 18332 44564 18460
rect 47395 18459 47453 18460
rect 46243 18416 46301 18417
rect 47404 18416 47444 18459
rect 47683 18416 47741 18417
rect 49516 18416 49556 18460
rect 51811 18459 51869 18460
rect 51331 18416 51389 18417
rect 44611 18376 44620 18416
rect 44660 18376 45484 18416
rect 45524 18376 45533 18416
rect 46158 18376 46252 18416
rect 46292 18376 46301 18416
rect 46819 18376 46828 18416
rect 46868 18376 47444 18416
rect 47491 18376 47500 18416
rect 47540 18376 47692 18416
rect 47732 18376 47741 18416
rect 48739 18376 48748 18416
rect 48788 18376 49556 18416
rect 51246 18376 51340 18416
rect 51380 18376 51389 18416
rect 46243 18375 46301 18376
rect 47683 18375 47741 18376
rect 51331 18375 51389 18376
rect 33283 18292 33292 18332
rect 33332 18292 35404 18332
rect 35444 18292 35453 18332
rect 44227 18292 44236 18332
rect 44276 18292 44564 18332
rect 45859 18292 45868 18332
rect 45908 18292 48460 18332
rect 48500 18292 49420 18332
rect 49460 18292 49469 18332
rect 49891 18292 49900 18332
rect 49940 18292 51724 18332
rect 51764 18292 51773 18332
rect 33283 18291 33341 18292
rect 33484 18248 33524 18292
rect 35395 18291 35453 18292
rect 40195 18248 40253 18249
rect 33475 18208 33484 18248
rect 33524 18208 33533 18248
rect 40110 18208 40204 18248
rect 40244 18208 40253 18248
rect 42883 18208 42892 18248
rect 42932 18208 46540 18248
rect 46580 18208 49324 18248
rect 49364 18208 49373 18248
rect 40195 18207 40253 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 3907 18124 3916 18164
rect 3956 18124 8620 18164
rect 8660 18124 8669 18164
rect 15103 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 15489 18164
rect 23011 18124 23020 18164
rect 23060 18124 24172 18164
rect 24212 18124 24221 18164
rect 26382 18124 26476 18164
rect 26516 18124 26525 18164
rect 27103 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 27489 18164
rect 28771 18124 28780 18164
rect 28820 18124 31756 18164
rect 31796 18124 31805 18164
rect 33100 18124 33580 18164
rect 33620 18124 33629 18164
rect 39103 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 39489 18164
rect 42019 18124 42028 18164
rect 42068 18124 45292 18164
rect 45332 18124 45964 18164
rect 46004 18124 48268 18164
rect 48308 18124 48317 18164
rect 50563 18124 50572 18164
rect 50612 18124 52780 18164
rect 52820 18124 52829 18164
rect 26467 18123 26525 18124
rect 28780 18080 28820 18124
rect 50572 18080 50612 18124
rect 3811 18040 3820 18080
rect 3860 18040 23596 18080
rect 23636 18040 23645 18080
rect 24547 18040 24556 18080
rect 24596 18040 25420 18080
rect 25460 18040 27916 18080
rect 27956 18040 28820 18080
rect 41539 18040 41548 18080
rect 41588 18040 43220 18080
rect 44707 18040 44716 18080
rect 44756 18040 44908 18080
rect 44948 18040 45676 18080
rect 45716 18040 50612 18080
rect 43180 17996 43220 18040
rect 8611 17956 8620 17996
rect 8660 17956 8908 17996
rect 8948 17956 8957 17996
rect 22435 17956 22444 17996
rect 22484 17956 22732 17996
rect 22772 17956 27436 17996
rect 27476 17956 30220 17996
rect 30260 17956 30269 17996
rect 41059 17956 41068 17996
rect 41108 17956 42028 17996
rect 42068 17956 42316 17996
rect 42356 17956 42365 17996
rect 43180 17956 45868 17996
rect 45908 17956 45917 17996
rect 46339 17956 46348 17996
rect 46388 17956 46732 17996
rect 46772 17956 46781 17996
rect 26467 17912 26525 17913
rect 22627 17872 22636 17912
rect 22676 17872 23348 17912
rect 24163 17872 24172 17912
rect 24212 17872 26420 17912
rect 1699 17788 1708 17828
rect 1748 17788 7948 17828
rect 7988 17788 9580 17828
rect 9620 17788 9629 17828
rect 23308 17744 23348 17872
rect 26380 17828 26420 17872
rect 26467 17872 26476 17912
rect 26516 17872 29740 17912
rect 29780 17872 29789 17912
rect 38563 17872 38572 17912
rect 38612 17872 48212 17912
rect 48451 17872 48460 17912
rect 48500 17872 48940 17912
rect 48980 17872 48989 17912
rect 49411 17872 49420 17912
rect 49460 17872 50572 17912
rect 50612 17872 50621 17912
rect 26467 17871 26525 17872
rect 26371 17788 26380 17828
rect 26420 17788 31276 17828
rect 31316 17788 31325 17828
rect 26467 17744 26525 17745
rect 38572 17744 38612 17872
rect 48172 17828 48212 17872
rect 42691 17788 42700 17828
rect 42740 17788 43948 17828
rect 43988 17788 43997 17828
rect 48172 17788 50476 17828
rect 50516 17788 50525 17828
rect 21667 17704 21676 17744
rect 21716 17704 22636 17744
rect 22676 17704 22685 17744
rect 22819 17704 22828 17744
rect 22868 17704 23212 17744
rect 23252 17704 23261 17744
rect 23308 17704 26476 17744
rect 26516 17704 26525 17744
rect 27715 17704 27724 17744
rect 27764 17704 27916 17744
rect 27956 17704 27965 17744
rect 31651 17704 31660 17744
rect 31700 17704 32236 17744
rect 32276 17704 32285 17744
rect 33283 17704 33292 17744
rect 33332 17704 34156 17744
rect 34196 17704 34205 17744
rect 36547 17704 36556 17744
rect 36596 17704 36844 17744
rect 36884 17704 38612 17744
rect 39811 17704 39820 17744
rect 39860 17704 41932 17744
rect 41972 17704 41981 17744
rect 42115 17704 42124 17744
rect 42164 17704 42892 17744
rect 42932 17704 44140 17744
rect 44180 17704 44189 17744
rect 50083 17704 50092 17744
rect 50132 17704 50380 17744
rect 50420 17704 51916 17744
rect 51956 17704 51965 17744
rect 5923 17620 5932 17660
rect 5972 17620 8044 17660
rect 8084 17620 8093 17660
rect 22636 17576 22676 17704
rect 26467 17703 26525 17704
rect 25507 17660 25565 17661
rect 22723 17620 22732 17660
rect 22772 17620 23116 17660
rect 23156 17620 23165 17660
rect 25422 17620 25516 17660
rect 25556 17620 25565 17660
rect 30019 17620 30028 17660
rect 30068 17620 30412 17660
rect 30452 17620 30461 17660
rect 42787 17620 42796 17660
rect 42836 17620 43180 17660
rect 43220 17620 43229 17660
rect 45955 17620 45964 17660
rect 46004 17620 46348 17660
rect 46388 17620 46397 17660
rect 25507 17619 25565 17620
rect 46723 17576 46781 17577
rect 22636 17536 26764 17576
rect 26804 17536 29932 17576
rect 29972 17536 31564 17576
rect 31604 17536 32524 17576
rect 32564 17536 32573 17576
rect 46147 17536 46156 17576
rect 46196 17536 46444 17576
rect 46484 17536 46732 17576
rect 46772 17536 48748 17576
rect 48788 17536 48797 17576
rect 46723 17535 46781 17536
rect 41059 17452 41068 17492
rect 41108 17452 41548 17492
rect 41588 17452 41597 17492
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 16343 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 16729 17408
rect 22531 17368 22540 17408
rect 22580 17368 22732 17408
rect 22772 17368 25516 17408
rect 25556 17368 25565 17408
rect 26851 17368 26860 17408
rect 26900 17368 26909 17408
rect 28343 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 28729 17408
rect 31939 17368 31948 17408
rect 31988 17368 33004 17408
rect 33044 17368 33292 17408
rect 33332 17368 33341 17408
rect 40343 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 40729 17408
rect 47971 17368 47980 17408
rect 48020 17368 48940 17408
rect 48980 17368 48989 17408
rect 0 17348 80 17368
rect 26860 17240 26900 17368
rect 32803 17324 32861 17325
rect 30508 17284 32812 17324
rect 32852 17284 32861 17324
rect 30508 17240 30548 17284
rect 32803 17283 32861 17284
rect 36844 17284 37132 17324
rect 37172 17284 37181 17324
rect 41059 17284 41068 17324
rect 41108 17284 43372 17324
rect 43412 17284 46828 17324
rect 46868 17284 46877 17324
rect 48835 17284 48844 17324
rect 48884 17284 49132 17324
rect 49172 17284 49181 17324
rect 51331 17284 51340 17324
rect 51380 17284 52012 17324
rect 52052 17284 52061 17324
rect 52387 17284 52396 17324
rect 52436 17284 54437 17324
rect 54477 17284 54486 17324
rect 36844 17240 36884 17284
rect 54307 17240 54365 17241
rect 55075 17240 55133 17241
rect 58243 17240 58301 17241
rect 75715 17240 75773 17241
rect 1699 17200 1708 17240
rect 1748 17200 2476 17240
rect 2516 17200 8812 17240
rect 8852 17200 8861 17240
rect 26860 17200 29164 17240
rect 29204 17200 29213 17240
rect 30468 17200 30508 17240
rect 30548 17200 30557 17240
rect 36163 17200 36172 17240
rect 36212 17200 36884 17240
rect 36931 17200 36940 17240
rect 36980 17200 37420 17240
rect 37460 17200 37469 17240
rect 48259 17200 48268 17240
rect 48308 17200 49228 17240
rect 49268 17200 49277 17240
rect 50659 17200 50668 17240
rect 50708 17200 51436 17240
rect 51476 17200 52684 17240
rect 52724 17200 53836 17240
rect 53876 17200 53885 17240
rect 54307 17200 54316 17240
rect 54385 17200 54451 17240
rect 54508 17200 54855 17240
rect 54895 17200 54904 17240
rect 55075 17200 55084 17240
rect 55124 17200 55145 17240
rect 55185 17200 55219 17240
rect 58243 17200 58252 17240
rect 58292 17200 58345 17240
rect 58385 17200 58394 17240
rect 61536 17200 61545 17240
rect 61585 17200 61804 17240
rect 61844 17200 61853 17240
rect 62336 17200 62345 17240
rect 62385 17200 62708 17240
rect 54307 17199 54365 17200
rect 40867 17156 40925 17157
rect 52291 17156 52349 17157
rect 54508 17156 54548 17200
rect 55075 17199 55133 17200
rect 58243 17199 58301 17200
rect 57859 17156 57917 17157
rect 40003 17116 40012 17156
rect 40052 17116 40876 17156
rect 40916 17116 40925 17156
rect 49891 17116 49900 17156
rect 49940 17116 51340 17156
rect 51380 17116 51389 17156
rect 52206 17116 52300 17156
rect 52340 17116 52349 17156
rect 52483 17116 52492 17156
rect 52532 17116 53655 17156
rect 53695 17116 53704 17156
rect 54028 17116 54055 17156
rect 54095 17116 54104 17156
rect 54499 17116 54508 17156
rect 54548 17116 54557 17156
rect 57859 17116 57868 17156
rect 57908 17116 57945 17156
rect 57985 17116 58003 17156
rect 40867 17115 40925 17116
rect 52291 17115 52349 17116
rect 52579 17072 52637 17073
rect 22915 17032 22924 17072
rect 22964 17032 24556 17072
rect 24596 17032 24605 17072
rect 26467 17032 26476 17072
rect 26516 17032 26860 17072
rect 26900 17032 26909 17072
rect 27043 17032 27052 17072
rect 27092 17032 27820 17072
rect 27860 17032 27869 17072
rect 30691 17032 30700 17072
rect 30740 17032 31948 17072
rect 31988 17032 31997 17072
rect 33955 17032 33964 17072
rect 34004 17032 34540 17072
rect 34580 17032 34589 17072
rect 38563 17032 38572 17072
rect 38612 17032 39724 17072
rect 39764 17032 39773 17072
rect 52195 17032 52204 17072
rect 52244 17032 52588 17072
rect 52628 17032 52637 17072
rect 52579 17031 52637 17032
rect 52771 17072 52829 17073
rect 52771 17032 52780 17072
rect 52820 17032 53932 17072
rect 53972 17032 53981 17072
rect 52771 17031 52829 17032
rect 46147 16988 46205 16989
rect 54028 16988 54068 17116
rect 57859 17115 57917 17116
rect 54691 17072 54749 17073
rect 62668 17072 62708 17200
rect 75715 17200 75724 17240
rect 75764 17200 75945 17240
rect 75985 17200 75994 17240
rect 75715 17199 75773 17200
rect 64579 17116 64588 17156
rect 64628 17116 64855 17156
rect 64895 17116 64904 17156
rect 66595 17116 66604 17156
rect 66644 17116 66855 17156
rect 66895 17116 66904 17156
rect 71395 17116 71404 17156
rect 71444 17116 71655 17156
rect 71695 17116 71704 17156
rect 78979 17116 78988 17156
rect 79028 17116 79372 17156
rect 79412 17116 79655 17156
rect 79695 17116 79704 17156
rect 54403 17032 54412 17072
rect 54452 17032 54700 17072
rect 54740 17032 54745 17072
rect 54785 17032 54835 17072
rect 62659 17032 62668 17072
rect 62708 17032 62717 17072
rect 54691 17031 54749 17032
rect 2659 16948 2668 16988
rect 2708 16948 5452 16988
rect 5492 16948 5501 16988
rect 41923 16948 41932 16988
rect 41972 16948 42124 16988
rect 42164 16948 42604 16988
rect 42644 16948 42653 16988
rect 45667 16948 45676 16988
rect 45716 16948 46156 16988
rect 46196 16948 48652 16988
rect 48692 16948 51476 16988
rect 52387 16948 52396 16988
rect 52436 16948 54068 16988
rect 46147 16947 46205 16948
rect 36643 16904 36701 16905
rect 51436 16904 51476 16948
rect 33964 16864 34348 16904
rect 34388 16864 36652 16904
rect 36692 16864 36701 16904
rect 37123 16864 37132 16904
rect 37172 16864 39764 16904
rect 40867 16864 40876 16904
rect 40916 16864 41356 16904
rect 41396 16864 41836 16904
rect 41876 16864 41885 16904
rect 42883 16864 42892 16904
rect 42932 16864 44044 16904
rect 44084 16864 44093 16904
rect 44707 16864 44716 16904
rect 44756 16864 45388 16904
rect 45428 16864 47212 16904
rect 47252 16864 48268 16904
rect 48308 16864 48317 16904
rect 49219 16864 49228 16904
rect 49268 16864 51340 16904
rect 51380 16864 51389 16904
rect 51436 16864 64684 16904
rect 64724 16864 64733 16904
rect 27523 16820 27581 16821
rect 29635 16820 29693 16821
rect 27427 16780 27436 16820
rect 27476 16780 27532 16820
rect 27572 16780 27581 16820
rect 29550 16780 29644 16820
rect 29684 16780 29693 16820
rect 27523 16779 27581 16780
rect 29635 16779 29693 16780
rect 33964 16736 34004 16864
rect 36643 16863 36701 16864
rect 39724 16821 39764 16864
rect 39715 16820 39773 16821
rect 49027 16820 49085 16821
rect 37027 16780 37036 16820
rect 37076 16780 37708 16820
rect 37748 16780 37757 16820
rect 39630 16780 39724 16820
rect 39764 16780 39773 16820
rect 41251 16780 41260 16820
rect 41300 16780 41740 16820
rect 41780 16780 41789 16820
rect 45091 16780 45100 16820
rect 45140 16780 45868 16820
rect 45908 16780 49036 16820
rect 49076 16780 49324 16820
rect 49364 16780 49373 16820
rect 49891 16780 49900 16820
rect 49940 16780 52204 16820
rect 52244 16780 52253 16820
rect 39715 16779 39773 16780
rect 49027 16779 49085 16780
rect 49900 16736 49940 16780
rect 33955 16696 33964 16736
rect 34004 16696 34013 16736
rect 43843 16696 43852 16736
rect 43892 16696 44524 16736
rect 44564 16696 49940 16736
rect 50467 16696 50476 16736
rect 50516 16696 55468 16736
rect 55508 16696 55517 16736
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 15103 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 15489 16652
rect 27103 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 27489 16652
rect 39103 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 39489 16652
rect 39907 16612 39916 16652
rect 39956 16612 42700 16652
rect 42740 16612 43220 16652
rect 50851 16612 50860 16652
rect 50900 16612 55660 16652
rect 55700 16612 55948 16652
rect 55988 16612 55997 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 43180 16484 43220 16612
rect 45955 16528 45964 16568
rect 46004 16528 46252 16568
rect 46292 16528 46301 16568
rect 53827 16528 53836 16568
rect 53876 16528 65356 16568
rect 65396 16528 65405 16568
rect 4195 16444 4204 16484
rect 4244 16444 4876 16484
rect 4916 16444 9388 16484
rect 9428 16444 9437 16484
rect 37315 16444 37324 16484
rect 37364 16444 37996 16484
rect 38036 16444 38045 16484
rect 43180 16444 57292 16484
rect 57332 16444 57341 16484
rect 61699 16444 61708 16484
rect 61748 16444 62188 16484
rect 62228 16444 62237 16484
rect 2371 16360 2380 16400
rect 2420 16360 4012 16400
rect 4052 16360 7660 16400
rect 7700 16360 7709 16400
rect 33475 16360 33484 16400
rect 33524 16360 33676 16400
rect 33716 16360 37420 16400
rect 37460 16360 37469 16400
rect 61699 16316 61757 16317
rect 33571 16276 33580 16316
rect 33620 16276 38036 16316
rect 61614 16276 61708 16316
rect 61748 16276 61757 16316
rect 27523 16232 27581 16233
rect 37996 16232 38036 16276
rect 61699 16275 61757 16276
rect 46243 16232 46301 16233
rect 52771 16232 52829 16233
rect 55075 16232 55133 16233
rect 58531 16232 58589 16233
rect 64963 16232 65021 16233
rect 70147 16232 70205 16233
rect 75715 16232 75773 16233
rect 77635 16232 77693 16233
rect 78883 16232 78941 16233
rect 5827 16192 5836 16232
rect 5876 16192 6316 16232
rect 6356 16192 7084 16232
rect 7124 16192 7133 16232
rect 27438 16192 27532 16232
rect 27572 16192 29644 16232
rect 29684 16192 29693 16232
rect 32515 16192 32524 16232
rect 32564 16192 34732 16232
rect 34772 16192 36268 16232
rect 36308 16192 36317 16232
rect 36451 16192 36460 16232
rect 36500 16192 37804 16232
rect 37844 16192 37853 16232
rect 37987 16192 37996 16232
rect 38036 16192 38045 16232
rect 39619 16192 39628 16232
rect 39668 16192 40108 16232
rect 40148 16192 40157 16232
rect 42499 16192 42508 16232
rect 42548 16192 42892 16232
rect 42932 16192 43220 16232
rect 46158 16192 46252 16232
rect 46292 16192 46301 16232
rect 48643 16192 48652 16232
rect 48692 16192 49420 16232
rect 49460 16192 49469 16232
rect 52686 16192 52780 16232
rect 52820 16192 52829 16232
rect 54787 16192 54796 16232
rect 54836 16192 55084 16232
rect 55124 16192 55133 16232
rect 56515 16192 56524 16232
rect 56564 16192 56573 16232
rect 58446 16192 58540 16232
rect 58580 16192 58589 16232
rect 60163 16192 60172 16232
rect 60212 16192 61900 16232
rect 61940 16192 62380 16232
rect 62420 16192 62429 16232
rect 64878 16192 64972 16232
rect 65012 16192 65021 16232
rect 66787 16192 66796 16232
rect 66836 16192 67372 16232
rect 67412 16192 67421 16232
rect 67939 16192 67948 16232
rect 67988 16192 69004 16232
rect 69044 16192 69053 16232
rect 70062 16192 70156 16232
rect 70196 16192 70205 16232
rect 74851 16192 74860 16232
rect 74900 16192 75340 16232
rect 75380 16192 75389 16232
rect 75630 16192 75724 16232
rect 75764 16192 75773 16232
rect 77155 16192 77164 16232
rect 77204 16192 77644 16232
rect 77684 16192 77693 16232
rect 78798 16192 78892 16232
rect 78932 16192 78941 16232
rect 27523 16191 27581 16192
rect 43180 16148 43220 16192
rect 46243 16191 46301 16192
rect 52771 16191 52829 16192
rect 55075 16191 55133 16192
rect 56524 16148 56564 16192
rect 58531 16191 58589 16192
rect 64963 16191 65021 16192
rect 70147 16191 70205 16192
rect 75715 16191 75773 16192
rect 77635 16191 77693 16192
rect 78883 16191 78941 16192
rect 2563 16108 2572 16148
rect 2612 16108 2956 16148
rect 2996 16108 21964 16148
rect 22004 16108 22013 16148
rect 27427 16108 27436 16148
rect 27476 16108 27820 16148
rect 27860 16108 27869 16148
rect 34915 16108 34924 16148
rect 34964 16108 35980 16148
rect 36020 16108 37036 16148
rect 37076 16108 37085 16148
rect 43180 16108 45580 16148
rect 45620 16108 56564 16148
rect 56620 16108 61556 16148
rect 61603 16108 61612 16148
rect 61652 16108 62668 16148
rect 62708 16108 62717 16148
rect 67267 16108 67276 16148
rect 67316 16108 69388 16148
rect 69428 16108 69437 16148
rect 71971 16108 71980 16148
rect 72020 16108 74956 16148
rect 74996 16108 75005 16148
rect 3619 16024 3628 16064
rect 3668 16024 6796 16064
rect 6836 16024 6845 16064
rect 6979 16024 6988 16064
rect 7028 16024 36172 16064
rect 36212 16024 36221 16064
rect 41635 16024 41644 16064
rect 41684 16024 44332 16064
rect 44372 16024 44524 16064
rect 44564 16024 44573 16064
rect 45475 16024 45484 16064
rect 45524 16024 56140 16064
rect 56180 16024 56189 16064
rect 51907 15980 51965 15981
rect 56620 15980 56660 16108
rect 61516 16064 61556 16108
rect 68515 16064 68573 16065
rect 57283 16024 57292 16064
rect 57332 16024 61132 16064
rect 61172 16024 61420 16064
rect 61460 16024 61469 16064
rect 61516 16024 63532 16064
rect 63572 16024 63581 16064
rect 68430 16024 68524 16064
rect 68564 16024 68573 16064
rect 68515 16023 68573 16024
rect 69091 16064 69149 16065
rect 77347 16064 77405 16065
rect 69091 16024 69100 16064
rect 69140 16024 70527 16064
rect 70567 16024 70576 16064
rect 76579 16024 76588 16064
rect 76628 16024 77356 16064
rect 77396 16024 77405 16064
rect 69091 16023 69149 16024
rect 77347 16023 77405 16024
rect 2179 15940 2188 15980
rect 2228 15940 2668 15980
rect 2708 15940 21580 15980
rect 21620 15940 21629 15980
rect 40003 15940 40012 15980
rect 40052 15940 40780 15980
rect 40820 15940 40829 15980
rect 51907 15940 51916 15980
rect 51956 15940 52012 15980
rect 52052 15940 52061 15980
rect 55459 15940 55468 15980
rect 55508 15940 56660 15980
rect 59491 15940 59500 15980
rect 59540 15940 66124 15980
rect 66164 15940 66173 15980
rect 69091 15940 69100 15980
rect 69140 15940 69772 15980
rect 69812 15940 69821 15980
rect 51907 15939 51965 15940
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 6787 15856 6796 15896
rect 6836 15856 8716 15896
rect 8756 15856 8765 15896
rect 16343 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 16729 15896
rect 28343 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 28729 15896
rect 33955 15856 33964 15896
rect 34004 15856 34636 15896
rect 34676 15856 34685 15896
rect 37411 15856 37420 15896
rect 37460 15856 40052 15896
rect 40343 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 40729 15896
rect 43267 15856 43276 15896
rect 43316 15856 45964 15896
rect 46004 15856 46013 15896
rect 49891 15856 49900 15896
rect 49940 15856 49949 15896
rect 51427 15856 51436 15896
rect 51476 15856 51820 15896
rect 51860 15856 52972 15896
rect 53012 15856 53021 15896
rect 53155 15856 53164 15896
rect 53204 15856 53452 15896
rect 53492 15856 53501 15896
rect 60652 15856 61804 15896
rect 61844 15856 62092 15896
rect 62132 15856 62141 15896
rect 40012 15812 40052 15856
rect 49900 15812 49940 15856
rect 60652 15813 60692 15856
rect 60643 15812 60701 15813
rect 29731 15772 29740 15812
rect 29780 15772 32908 15812
rect 32948 15772 33484 15812
rect 33524 15772 36172 15812
rect 36212 15772 36221 15812
rect 40003 15772 40012 15812
rect 40052 15772 40061 15812
rect 49900 15772 51628 15812
rect 51668 15772 52012 15812
rect 52052 15772 52061 15812
rect 54595 15772 54604 15812
rect 54644 15772 58924 15812
rect 58964 15772 58973 15812
rect 60643 15772 60652 15812
rect 60692 15772 60701 15812
rect 76963 15772 76972 15812
rect 77012 15772 78412 15812
rect 78452 15772 78461 15812
rect 60643 15771 60701 15772
rect 0 15728 80 15748
rect 47683 15728 47741 15729
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 2179 15688 2188 15728
rect 2228 15688 3436 15728
rect 3476 15688 4300 15728
rect 4340 15688 4349 15728
rect 30979 15688 30988 15728
rect 31028 15688 33868 15728
rect 33908 15688 33917 15728
rect 45475 15688 45484 15728
rect 45524 15688 47692 15728
rect 47732 15688 47741 15728
rect 52771 15688 52780 15728
rect 52820 15688 53164 15728
rect 53204 15688 53213 15728
rect 64483 15688 64492 15728
rect 64532 15688 64780 15728
rect 64820 15688 67852 15728
rect 67892 15688 72556 15728
rect 72596 15688 72605 15728
rect 0 15668 80 15688
rect 47683 15687 47741 15688
rect 33091 15644 33149 15645
rect 32323 15604 32332 15644
rect 32372 15604 32812 15644
rect 32852 15604 33100 15644
rect 33140 15604 33149 15644
rect 33091 15603 33149 15604
rect 33196 15604 34636 15644
rect 34676 15604 34685 15644
rect 39619 15604 39628 15644
rect 39668 15604 42028 15644
rect 42068 15604 42220 15644
rect 42260 15604 43084 15644
rect 43124 15604 43133 15644
rect 45571 15604 45580 15644
rect 45620 15604 46252 15644
rect 46292 15604 47404 15644
rect 47444 15604 48076 15644
rect 48116 15604 48125 15644
rect 49123 15604 49132 15644
rect 49172 15604 51148 15644
rect 51188 15604 53644 15644
rect 53684 15604 53693 15644
rect 33196 15560 33236 15604
rect 47971 15560 48029 15561
rect 4195 15520 4204 15560
rect 4244 15520 4780 15560
rect 4820 15520 4829 15560
rect 31939 15520 31948 15560
rect 31988 15520 33004 15560
rect 33044 15520 33236 15560
rect 34435 15520 34444 15560
rect 34484 15520 34493 15560
rect 36067 15520 36076 15560
rect 36116 15520 36844 15560
rect 36884 15520 36893 15560
rect 37507 15520 37516 15560
rect 37556 15520 37565 15560
rect 39139 15520 39148 15560
rect 39188 15520 40204 15560
rect 40244 15520 40588 15560
rect 40628 15520 40637 15560
rect 46051 15520 46060 15560
rect 46100 15520 46444 15560
rect 46484 15520 46493 15560
rect 47886 15520 47980 15560
rect 48020 15520 48029 15560
rect 49987 15520 49996 15560
rect 50036 15520 50764 15560
rect 50804 15520 51052 15560
rect 51092 15520 51101 15560
rect 51811 15520 51820 15560
rect 51860 15520 52588 15560
rect 52628 15520 53204 15560
rect 61987 15520 61996 15560
rect 62036 15520 64972 15560
rect 65012 15520 65021 15560
rect 70723 15520 70732 15560
rect 70772 15520 75148 15560
rect 75188 15520 75197 15560
rect 835 15436 844 15476
rect 884 15436 4684 15476
rect 4724 15436 6988 15476
rect 7028 15436 7037 15476
rect 29827 15436 29836 15476
rect 29876 15436 33388 15476
rect 33428 15436 33437 15476
rect 2860 15140 2900 15436
rect 4771 15392 4829 15393
rect 4483 15352 4492 15392
rect 4532 15352 4780 15392
rect 4820 15352 9004 15392
rect 9044 15352 9053 15392
rect 4771 15351 4829 15352
rect 33004 15308 33044 15436
rect 33187 15392 33245 15393
rect 34444 15392 34484 15520
rect 37516 15476 37556 15520
rect 47971 15519 48029 15520
rect 53164 15476 53204 15520
rect 36259 15436 36268 15476
rect 36308 15436 37556 15476
rect 53155 15436 53164 15476
rect 53204 15436 53213 15476
rect 55555 15436 55564 15476
rect 55604 15436 63284 15476
rect 62947 15392 63005 15393
rect 33187 15352 33196 15392
rect 33236 15352 35116 15392
rect 35156 15352 35165 15392
rect 39235 15352 39244 15392
rect 39284 15352 43660 15392
rect 43700 15352 44236 15392
rect 44276 15352 44285 15392
rect 47203 15352 47212 15392
rect 47252 15352 47788 15392
rect 47828 15352 50380 15392
rect 50420 15352 62956 15392
rect 62996 15352 63005 15392
rect 33187 15351 33245 15352
rect 62947 15351 63005 15352
rect 63244 15308 63284 15436
rect 63331 15392 63389 15393
rect 64972 15392 65012 15520
rect 66211 15436 66220 15476
rect 66260 15436 68716 15476
rect 68756 15436 74284 15476
rect 74324 15436 74333 15476
rect 63331 15352 63340 15392
rect 63380 15352 64108 15392
rect 64148 15352 64157 15392
rect 64972 15352 69812 15392
rect 69859 15352 69868 15392
rect 69908 15352 74668 15392
rect 74708 15352 74717 15392
rect 63331 15351 63389 15352
rect 69772 15308 69812 15352
rect 2947 15268 2956 15308
rect 2996 15268 3436 15308
rect 3476 15268 3485 15308
rect 31747 15268 31756 15308
rect 31796 15268 32044 15308
rect 32084 15268 32093 15308
rect 32995 15268 33004 15308
rect 33044 15268 33053 15308
rect 48931 15268 48940 15308
rect 48980 15268 49996 15308
rect 50036 15268 50045 15308
rect 52483 15268 52492 15308
rect 52532 15268 53356 15308
rect 53396 15268 55564 15308
rect 55604 15268 55613 15308
rect 56995 15268 57004 15308
rect 57044 15268 61612 15308
rect 61652 15268 61661 15308
rect 62371 15268 62380 15308
rect 62420 15268 62956 15308
rect 62996 15268 63005 15308
rect 63244 15268 65740 15308
rect 65780 15268 65789 15308
rect 69772 15268 70540 15308
rect 70580 15268 71116 15308
rect 71156 15268 71165 15308
rect 73795 15268 73804 15308
rect 73844 15268 75244 15308
rect 75284 15268 75628 15308
rect 75668 15268 75677 15308
rect 62956 15224 62996 15268
rect 7459 15184 7468 15224
rect 7508 15184 45196 15224
rect 45236 15184 45245 15224
rect 62956 15184 72172 15224
rect 72212 15184 72221 15224
rect 2851 15100 2860 15140
rect 2900 15100 2909 15140
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 15103 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 15489 15140
rect 27103 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 27489 15140
rect 39103 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 39489 15140
rect 51103 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 51489 15140
rect 63103 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 63489 15140
rect 70819 15100 70828 15140
rect 70868 15100 71308 15140
rect 71348 15100 71357 15140
rect 75103 15100 75112 15140
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75480 15100 75489 15140
rect 60739 15056 60797 15057
rect 60739 15016 60748 15056
rect 60788 15016 69868 15056
rect 69908 15016 69917 15056
rect 60739 15015 60797 15016
rect 1027 14932 1036 14972
rect 1076 14932 1996 14972
rect 2036 14932 2045 14972
rect 38179 14932 38188 14972
rect 38228 14932 39436 14972
rect 39476 14932 39485 14972
rect 45571 14932 45580 14972
rect 45620 14932 46156 14972
rect 46196 14932 46205 14972
rect 61612 14932 70636 14972
rect 70676 14932 70685 14972
rect 78595 14932 78604 14972
rect 78644 14932 79180 14972
rect 79220 14932 79229 14972
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 1795 14848 1804 14888
rect 1844 14848 2764 14888
rect 2804 14848 2813 14888
rect 35587 14848 35596 14888
rect 35636 14848 36940 14888
rect 36980 14848 36989 14888
rect 57187 14848 57196 14888
rect 57236 14848 57484 14888
rect 57524 14848 57533 14888
rect 0 14828 80 14848
rect 46723 14804 46781 14805
rect 47971 14804 48029 14805
rect 32995 14764 33004 14804
rect 33044 14764 35500 14804
rect 35540 14764 36076 14804
rect 36116 14764 36125 14804
rect 45763 14764 45772 14804
rect 45812 14764 46732 14804
rect 46772 14764 47980 14804
rect 48020 14764 48029 14804
rect 46723 14763 46781 14764
rect 47971 14763 48029 14764
rect 50755 14804 50813 14805
rect 61612 14804 61652 14932
rect 61891 14888 61949 14889
rect 61891 14848 61900 14888
rect 61940 14848 62764 14888
rect 62804 14848 70732 14888
rect 70772 14848 70781 14888
rect 73603 14848 73612 14888
rect 73652 14848 74092 14888
rect 74132 14848 74141 14888
rect 75619 14848 75628 14888
rect 75668 14848 75677 14888
rect 61891 14847 61949 14848
rect 67171 14804 67229 14805
rect 75628 14804 75668 14848
rect 50755 14764 50764 14804
rect 50804 14764 61612 14804
rect 61652 14764 61661 14804
rect 67086 14764 67180 14804
rect 67220 14764 74764 14804
rect 74804 14764 74813 14804
rect 75628 14764 75860 14804
rect 50755 14763 50813 14764
rect 67171 14763 67229 14764
rect 60739 14720 60797 14721
rect 75820 14720 75860 14764
rect 1507 14680 1516 14720
rect 1556 14680 2956 14720
rect 2996 14680 3005 14720
rect 5251 14680 5260 14720
rect 5300 14680 7468 14720
rect 7508 14680 7517 14720
rect 31171 14680 31180 14720
rect 31220 14680 34252 14720
rect 34292 14680 35212 14720
rect 35252 14680 36844 14720
rect 36884 14680 38092 14720
rect 38132 14680 38572 14720
rect 38612 14680 38621 14720
rect 41443 14680 41452 14720
rect 41492 14680 41501 14720
rect 42019 14680 42028 14720
rect 42068 14680 42604 14720
rect 42644 14680 42796 14720
rect 42836 14680 42845 14720
rect 43075 14680 43084 14720
rect 43124 14680 43372 14720
rect 43412 14680 43421 14720
rect 45859 14680 45868 14720
rect 45908 14680 46348 14720
rect 46388 14680 47308 14720
rect 47348 14680 47357 14720
rect 52291 14680 52300 14720
rect 52340 14680 56044 14720
rect 56084 14680 56093 14720
rect 56323 14680 56332 14720
rect 56372 14680 57580 14720
rect 57620 14680 59500 14720
rect 59540 14680 59549 14720
rect 60654 14680 60748 14720
rect 60788 14680 60797 14720
rect 61219 14680 61228 14720
rect 61268 14680 62284 14720
rect 62324 14680 62333 14720
rect 63811 14680 63820 14720
rect 63860 14680 64684 14720
rect 64724 14680 65164 14720
rect 65204 14680 65213 14720
rect 70627 14680 70636 14720
rect 70676 14680 75628 14720
rect 75668 14680 75677 14720
rect 75811 14680 75820 14720
rect 75860 14680 75869 14720
rect 4771 14596 4780 14636
rect 4820 14596 5164 14636
rect 5204 14596 5213 14636
rect 29923 14596 29932 14636
rect 29972 14596 31372 14636
rect 31412 14596 31421 14636
rect 39619 14596 39628 14636
rect 39668 14596 39677 14636
rect 32323 14552 32381 14553
rect 32131 14512 32140 14552
rect 32180 14512 32332 14552
rect 32372 14512 32381 14552
rect 39628 14552 39668 14596
rect 39628 14512 40012 14552
rect 40052 14512 40061 14552
rect 32323 14511 32381 14512
rect 4867 14468 4925 14469
rect 2947 14428 2956 14468
rect 2996 14428 4876 14468
rect 4916 14428 4925 14468
rect 41347 14428 41356 14468
rect 41396 14428 41405 14468
rect 4867 14427 4925 14428
rect 41356 14384 41396 14428
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 16343 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 16729 14384
rect 28343 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 28729 14384
rect 40343 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 40729 14384
rect 41059 14344 41068 14384
rect 41108 14344 41396 14384
rect 41452 14300 41492 14680
rect 49315 14636 49373 14637
rect 56044 14636 56084 14680
rect 60739 14679 60797 14680
rect 46243 14596 46252 14636
rect 46292 14596 49228 14636
rect 49268 14596 49324 14636
rect 49364 14596 49392 14636
rect 56044 14596 57676 14636
rect 57716 14596 57725 14636
rect 67555 14596 67564 14636
rect 67604 14596 68236 14636
rect 68276 14596 68285 14636
rect 74371 14596 74380 14636
rect 74420 14596 75052 14636
rect 75092 14596 75101 14636
rect 49315 14595 49373 14596
rect 46915 14512 46924 14552
rect 46964 14512 48364 14552
rect 48404 14512 48413 14552
rect 52675 14512 52684 14552
rect 52724 14512 56908 14552
rect 56948 14512 58828 14552
rect 58868 14512 58877 14552
rect 59491 14512 59500 14552
rect 59540 14512 61804 14552
rect 61844 14512 62188 14552
rect 62228 14512 63916 14552
rect 63956 14512 63965 14552
rect 70531 14512 70540 14552
rect 70580 14512 70828 14552
rect 70868 14512 70877 14552
rect 72163 14512 72172 14552
rect 72212 14512 73708 14552
rect 73748 14512 73757 14552
rect 74947 14512 74956 14552
rect 74996 14512 76012 14552
rect 76052 14512 78604 14552
rect 78644 14512 78653 14552
rect 52099 14428 52108 14468
rect 52148 14428 54412 14468
rect 54452 14428 55084 14468
rect 55124 14428 55948 14468
rect 55988 14428 58348 14468
rect 58388 14428 58397 14468
rect 62563 14428 62572 14468
rect 62612 14428 62621 14468
rect 70147 14428 70156 14468
rect 70196 14428 71020 14468
rect 71060 14428 71069 14468
rect 73603 14428 73612 14468
rect 73652 14428 74860 14468
rect 74900 14428 74909 14468
rect 58348 14384 58388 14428
rect 62572 14384 62612 14428
rect 46051 14344 46060 14384
rect 46100 14344 46540 14384
rect 46580 14344 47404 14384
rect 47444 14344 48652 14384
rect 48692 14344 48701 14384
rect 50563 14344 50572 14384
rect 50612 14344 51628 14384
rect 51668 14344 51677 14384
rect 52343 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 52729 14384
rect 58348 14344 59404 14384
rect 59444 14344 60460 14384
rect 60500 14344 61708 14384
rect 61748 14344 62476 14384
rect 62516 14344 62525 14384
rect 62572 14344 63724 14384
rect 63764 14344 63773 14384
rect 64343 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 64729 14384
rect 68323 14344 68332 14384
rect 68372 14344 68524 14384
rect 68564 14344 68573 14384
rect 69187 14344 69196 14384
rect 69236 14344 74188 14384
rect 74228 14344 74237 14384
rect 74371 14344 74380 14384
rect 74420 14344 74429 14384
rect 76343 14344 76352 14384
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76720 14344 76729 14384
rect 1603 14260 1612 14300
rect 1652 14260 2188 14300
rect 2228 14260 2380 14300
rect 2420 14260 3916 14300
rect 3956 14260 3965 14300
rect 39331 14260 39340 14300
rect 39380 14260 41164 14300
rect 41204 14260 41356 14300
rect 41396 14260 41492 14300
rect 57955 14260 57964 14300
rect 58004 14260 60652 14300
rect 60692 14260 66508 14300
rect 66548 14260 66557 14300
rect 66979 14260 66988 14300
rect 67028 14260 69100 14300
rect 69140 14260 69149 14300
rect 2275 14176 2284 14216
rect 2324 14176 2860 14216
rect 2900 14176 2909 14216
rect 32227 14176 32236 14216
rect 32276 14176 32716 14216
rect 32756 14176 32765 14216
rect 32995 14176 33004 14216
rect 33044 14176 34828 14216
rect 34868 14176 35404 14216
rect 35444 14176 35453 14216
rect 37795 14176 37804 14216
rect 37844 14176 38380 14216
rect 38420 14176 38429 14216
rect 39811 14176 39820 14216
rect 39860 14176 41260 14216
rect 41300 14176 42604 14216
rect 42644 14176 43220 14216
rect 50755 14176 50764 14216
rect 50804 14176 51340 14216
rect 51380 14176 51389 14216
rect 52195 14176 52204 14216
rect 52244 14176 73460 14216
rect 33004 14132 33044 14176
rect 43180 14132 43220 14176
rect 52771 14132 52829 14133
rect 4291 14092 4300 14132
rect 4340 14092 5260 14132
rect 5300 14092 5309 14132
rect 32323 14092 32332 14132
rect 32372 14092 33044 14132
rect 37411 14092 37420 14132
rect 37460 14092 38572 14132
rect 38612 14092 39148 14132
rect 39188 14092 39197 14132
rect 43171 14092 43180 14132
rect 43220 14092 43229 14132
rect 43363 14092 43372 14132
rect 43412 14092 43564 14132
rect 43604 14092 43613 14132
rect 44323 14092 44332 14132
rect 44372 14092 45868 14132
rect 45908 14092 46252 14132
rect 46292 14092 46301 14132
rect 47587 14092 47596 14132
rect 47636 14092 49036 14132
rect 49076 14092 49324 14132
rect 49364 14092 49373 14132
rect 51235 14092 51244 14132
rect 51284 14092 52780 14132
rect 52820 14092 52972 14132
rect 53012 14092 53021 14132
rect 61411 14092 61420 14132
rect 61460 14092 62380 14132
rect 62420 14092 62429 14132
rect 68803 14092 68812 14132
rect 68852 14092 69388 14132
rect 69428 14092 70060 14132
rect 70100 14092 70109 14132
rect 52771 14091 52829 14092
rect 0 14048 80 14068
rect 1987 14048 2045 14049
rect 57763 14048 57821 14049
rect 73420 14048 73460 14176
rect 74380 14048 74420 14344
rect 77155 14176 77164 14216
rect 77204 14176 78700 14216
rect 78740 14176 79372 14216
rect 79412 14176 79421 14216
rect 0 14008 1036 14048
rect 1076 14008 1085 14048
rect 1987 14008 1996 14048
rect 2036 14008 3052 14048
rect 3092 14008 4396 14048
rect 4436 14008 4445 14048
rect 31843 14008 31852 14048
rect 31892 14008 37228 14048
rect 37268 14008 37804 14048
rect 37844 14008 46156 14048
rect 46196 14008 46205 14048
rect 46531 14008 46540 14048
rect 46580 14008 47500 14048
rect 47540 14008 47788 14048
rect 47828 14008 47837 14048
rect 53827 14008 53836 14048
rect 53876 14008 54700 14048
rect 54740 14008 54749 14048
rect 57678 14008 57772 14048
rect 57812 14008 57821 14048
rect 60835 14008 60844 14048
rect 60884 14008 61844 14048
rect 62467 14008 62476 14048
rect 62516 14008 65932 14048
rect 65972 14008 66700 14048
rect 66740 14008 66749 14048
rect 69955 14008 69964 14048
rect 70004 14008 71116 14048
rect 71156 14008 72748 14048
rect 72788 14008 72797 14048
rect 73420 14008 74668 14048
rect 74708 14008 74717 14048
rect 77635 14008 77644 14048
rect 77684 14008 78220 14048
rect 78260 14008 78269 14048
rect 0 13988 80 14008
rect 1987 14007 2045 14008
rect 57763 14007 57821 14008
rect 61804 13964 61844 14008
rect 63907 13964 63965 13965
rect 1315 13924 1324 13964
rect 1364 13924 4300 13964
rect 4340 13924 4349 13964
rect 38467 13924 38476 13964
rect 38516 13924 38860 13964
rect 38900 13924 38909 13964
rect 39235 13924 39244 13964
rect 39284 13924 41068 13964
rect 41108 13924 41117 13964
rect 60547 13924 60556 13964
rect 60596 13924 61708 13964
rect 61748 13924 61757 13964
rect 61804 13924 62572 13964
rect 62612 13924 62621 13964
rect 63822 13924 63916 13964
rect 63956 13924 63965 13964
rect 64387 13924 64396 13964
rect 64436 13924 67084 13964
rect 67124 13924 67276 13964
rect 67316 13924 67325 13964
rect 68131 13924 68140 13964
rect 68180 13924 69868 13964
rect 69908 13924 69917 13964
rect 74947 13924 74956 13964
rect 74996 13924 75005 13964
rect 63907 13923 63965 13924
rect 69187 13880 69245 13881
rect 74956 13880 74996 13924
rect 36163 13840 36172 13880
rect 36212 13840 37324 13880
rect 37364 13840 38092 13880
rect 38132 13840 38141 13880
rect 40099 13840 40108 13880
rect 40148 13840 41932 13880
rect 41972 13840 42316 13880
rect 42356 13840 42365 13880
rect 53059 13840 53068 13880
rect 53108 13840 56428 13880
rect 56468 13840 58348 13880
rect 58388 13840 58397 13880
rect 65539 13840 65548 13880
rect 65588 13840 67372 13880
rect 67412 13840 67421 13880
rect 67555 13840 67564 13880
rect 67604 13840 68044 13880
rect 68084 13840 68093 13880
rect 69102 13840 69196 13880
rect 69236 13840 69245 13880
rect 69187 13839 69245 13840
rect 69292 13840 70924 13880
rect 70964 13840 74860 13880
rect 74900 13840 74996 13880
rect 68515 13796 68573 13797
rect 69292 13796 69332 13840
rect 739 13756 748 13796
rect 788 13756 1516 13796
rect 1556 13756 1565 13796
rect 4675 13756 4684 13796
rect 4724 13756 6604 13796
rect 6644 13756 6653 13796
rect 57859 13756 57868 13796
rect 57908 13756 59020 13796
rect 59060 13756 59069 13796
rect 68131 13756 68140 13796
rect 68180 13756 68524 13796
rect 68564 13756 68573 13796
rect 69283 13756 69292 13796
rect 69332 13756 69341 13796
rect 70819 13756 70828 13796
rect 70868 13756 75820 13796
rect 75860 13756 75869 13796
rect 68515 13755 68573 13756
rect 43459 13672 43468 13712
rect 43508 13672 43852 13712
rect 43892 13672 43901 13712
rect 54499 13672 54508 13712
rect 54548 13672 56524 13712
rect 56564 13672 57100 13712
rect 57140 13672 57149 13712
rect 67843 13672 67852 13712
rect 67892 13672 68044 13712
rect 68084 13672 68093 13712
rect 73891 13672 73900 13712
rect 73940 13672 74764 13712
rect 74804 13672 74813 13712
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 15103 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 15489 13628
rect 27103 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 27489 13628
rect 39103 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 39489 13628
rect 51103 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 51489 13628
rect 53539 13588 53548 13628
rect 53588 13588 56236 13628
rect 56276 13588 56285 13628
rect 63103 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 63489 13628
rect 68515 13588 68524 13628
rect 68564 13588 68716 13628
rect 68756 13588 69100 13628
rect 69140 13588 69149 13628
rect 75103 13588 75112 13628
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75480 13588 75489 13628
rect 2371 13504 2380 13544
rect 2420 13504 2764 13544
rect 2804 13504 2813 13544
rect 32707 13504 32716 13544
rect 32756 13504 37132 13544
rect 37172 13504 37181 13544
rect 47500 13504 56812 13544
rect 56852 13504 56861 13544
rect 57388 13504 57964 13544
rect 58004 13504 58013 13544
rect 69859 13504 69868 13544
rect 69908 13504 70156 13544
rect 70196 13504 70205 13544
rect 74851 13504 74860 13544
rect 74900 13504 75188 13544
rect 36643 13460 36701 13461
rect 47500 13460 47540 13504
rect 31651 13420 31660 13460
rect 31700 13420 32428 13460
rect 32468 13420 32812 13460
rect 32852 13420 32861 13460
rect 36259 13420 36268 13460
rect 36308 13420 36652 13460
rect 36692 13420 36701 13460
rect 40291 13420 40300 13460
rect 40340 13420 41548 13460
rect 41588 13420 41597 13460
rect 43267 13420 43276 13460
rect 43316 13420 45484 13460
rect 45524 13420 47540 13460
rect 47683 13460 47741 13461
rect 57388 13460 57428 13504
rect 74851 13460 74909 13461
rect 75148 13460 75188 13504
rect 47683 13420 47692 13460
rect 47732 13420 48076 13460
rect 48116 13420 48125 13460
rect 50851 13420 50860 13460
rect 50900 13420 51532 13460
rect 51572 13420 53452 13460
rect 53492 13420 56140 13460
rect 56180 13420 57388 13460
rect 57428 13420 57437 13460
rect 57484 13420 63532 13460
rect 63572 13420 63581 13460
rect 68419 13420 68428 13460
rect 68468 13420 68812 13460
rect 68852 13420 74860 13460
rect 74900 13420 74909 13460
rect 75139 13420 75148 13460
rect 75188 13420 75197 13460
rect 36643 13419 36701 13420
rect 47683 13419 47741 13420
rect 57484 13376 57524 13420
rect 74851 13419 74909 13420
rect 2467 13336 2476 13376
rect 2516 13336 2764 13376
rect 2804 13336 3340 13376
rect 3380 13336 3389 13376
rect 5443 13336 5452 13376
rect 5492 13336 6220 13376
rect 6260 13336 6269 13376
rect 42595 13336 42604 13376
rect 42644 13336 46060 13376
rect 46100 13336 46109 13376
rect 46540 13336 48460 13376
rect 48500 13336 48509 13376
rect 51811 13336 51820 13376
rect 51860 13336 57524 13376
rect 61603 13336 61612 13376
rect 61652 13336 62476 13376
rect 62516 13336 62525 13376
rect 64099 13336 64108 13376
rect 64148 13336 64396 13376
rect 64436 13336 64445 13376
rect 73420 13336 74380 13376
rect 74420 13336 74429 13376
rect 74563 13336 74572 13376
rect 74612 13336 74956 13376
rect 74996 13336 75092 13376
rect 2860 13252 4876 13292
rect 4916 13252 6700 13292
rect 6740 13252 6749 13292
rect 35395 13252 35404 13292
rect 35444 13252 36076 13292
rect 36116 13252 36125 13292
rect 36259 13252 36268 13292
rect 36308 13252 36596 13292
rect 0 13208 80 13228
rect 2860 13208 2900 13252
rect 36556 13208 36596 13252
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 1699 13168 1708 13208
rect 1748 13168 2900 13208
rect 5155 13168 5164 13208
rect 5204 13168 31852 13208
rect 31892 13168 31901 13208
rect 36547 13168 36556 13208
rect 36596 13168 37036 13208
rect 37076 13168 38860 13208
rect 38900 13168 38909 13208
rect 41731 13168 41740 13208
rect 41780 13168 42796 13208
rect 42836 13168 42845 13208
rect 0 13148 80 13168
rect 46540 13124 46580 13336
rect 47971 13292 48029 13293
rect 47491 13252 47500 13292
rect 47540 13252 47980 13292
rect 48020 13252 49516 13292
rect 49556 13252 49565 13292
rect 51619 13252 51628 13292
rect 51668 13252 55180 13292
rect 55220 13252 56908 13292
rect 56948 13252 56957 13292
rect 61987 13252 61996 13292
rect 62036 13252 62860 13292
rect 62900 13252 62909 13292
rect 67459 13252 67468 13292
rect 67508 13252 69100 13292
rect 69140 13252 69149 13292
rect 47971 13251 48029 13252
rect 49315 13208 49373 13209
rect 73420 13208 73460 13336
rect 75052 13208 75092 13336
rect 75715 13252 75724 13292
rect 75764 13252 77164 13292
rect 77204 13252 77213 13292
rect 76195 13208 76253 13209
rect 49315 13168 49324 13208
rect 49364 13168 50668 13208
rect 50708 13168 53260 13208
rect 53300 13168 53309 13208
rect 55363 13168 55372 13208
rect 55412 13168 56044 13208
rect 56084 13168 56093 13208
rect 56323 13168 56332 13208
rect 56372 13168 56660 13208
rect 56707 13168 56716 13208
rect 56756 13168 58540 13208
rect 58580 13168 58924 13208
rect 58964 13168 58973 13208
rect 61315 13168 61324 13208
rect 61364 13168 62284 13208
rect 62324 13168 63628 13208
rect 63668 13168 63677 13208
rect 63907 13168 63916 13208
rect 63956 13168 63965 13208
rect 68899 13168 68908 13208
rect 68948 13168 69580 13208
rect 69620 13168 69629 13208
rect 72163 13168 72172 13208
rect 72212 13168 73460 13208
rect 74275 13168 74284 13208
rect 74324 13168 74764 13208
rect 74804 13168 74813 13208
rect 75043 13168 75052 13208
rect 75092 13168 75820 13208
rect 75860 13168 75869 13208
rect 76195 13168 76204 13208
rect 76244 13168 76492 13208
rect 76532 13168 76541 13208
rect 49315 13167 49373 13168
rect 56620 13124 56660 13168
rect 63916 13124 63956 13168
rect 76195 13167 76253 13168
rect 3331 13084 3340 13124
rect 3380 13084 5356 13124
rect 5396 13084 5405 13124
rect 36835 13084 36844 13124
rect 36884 13084 39340 13124
rect 39380 13084 46580 13124
rect 49123 13084 49132 13124
rect 49172 13084 49420 13124
rect 49460 13084 49469 13124
rect 51715 13084 51724 13124
rect 51764 13084 55276 13124
rect 55316 13084 56428 13124
rect 56468 13084 56477 13124
rect 56620 13084 57716 13124
rect 62851 13084 62860 13124
rect 62900 13084 63956 13124
rect 74851 13124 74909 13125
rect 74851 13084 74860 13124
rect 74900 13084 74956 13124
rect 74996 13084 75005 13124
rect 75139 13084 75148 13124
rect 75188 13084 76972 13124
rect 77012 13084 77021 13124
rect 36355 13040 36413 13041
rect 57676 13040 57716 13084
rect 74851 13083 74909 13084
rect 57859 13040 57917 13041
rect 68899 13040 68957 13041
rect 1411 13000 1420 13040
rect 1460 13000 3628 13040
rect 3668 13000 3677 13040
rect 35107 13000 35116 13040
rect 35156 13000 36364 13040
rect 36404 13000 38284 13040
rect 38324 13000 38333 13040
rect 42691 13000 42700 13040
rect 42740 13000 43660 13040
rect 43700 13000 44428 13040
rect 44468 13000 44477 13040
rect 46243 13000 46252 13040
rect 46292 13000 46636 13040
rect 46676 13000 46685 13040
rect 48451 13000 48460 13040
rect 48500 13000 54604 13040
rect 54644 13000 54653 13040
rect 54883 13000 54892 13040
rect 54932 13000 56620 13040
rect 56660 13000 56669 13040
rect 57667 13000 57676 13040
rect 57716 13000 57725 13040
rect 57859 13000 57868 13040
rect 57908 13000 58002 13040
rect 61123 13000 61132 13040
rect 61172 13000 61996 13040
rect 62036 13000 62045 13040
rect 63811 13000 63820 13040
rect 63860 13000 64588 13040
rect 64628 13000 64637 13040
rect 68611 13000 68620 13040
rect 68660 13000 68908 13040
rect 68948 13000 68957 13040
rect 69475 13000 69484 13040
rect 69524 13000 70156 13040
rect 70196 13000 75532 13040
rect 75572 13000 75581 13040
rect 36355 12999 36413 13000
rect 57859 12999 57917 13000
rect 68899 12999 68957 13000
rect 62179 12916 62188 12956
rect 62228 12916 63532 12956
rect 63572 12916 64012 12956
rect 64052 12916 64061 12956
rect 68620 12916 69004 12956
rect 69044 12916 71596 12956
rect 71636 12916 73036 12956
rect 73076 12916 73420 12956
rect 73460 12916 73708 12956
rect 73748 12916 77644 12956
rect 77684 12916 77693 12956
rect 51907 12872 51965 12873
rect 68620 12872 68660 12916
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 16343 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 16729 12872
rect 28343 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 28729 12872
rect 40343 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 40729 12872
rect 42307 12832 42316 12872
rect 42356 12832 42988 12872
rect 43028 12832 47500 12872
rect 47540 12832 47549 12872
rect 49699 12832 49708 12872
rect 49748 12832 50380 12872
rect 50420 12832 50429 12872
rect 51822 12832 51916 12872
rect 51956 12832 51965 12872
rect 52343 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 52729 12872
rect 64343 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 64729 12872
rect 68611 12832 68620 12872
rect 68660 12832 68669 12872
rect 69763 12832 69772 12872
rect 69812 12832 70060 12872
rect 70100 12832 70109 12872
rect 76343 12832 76352 12872
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76720 12832 76729 12872
rect 51907 12831 51965 12832
rect 48451 12748 48460 12788
rect 48500 12748 49748 12788
rect 49708 12704 49748 12748
rect 53260 12748 59308 12788
rect 59348 12748 59357 12788
rect 67171 12748 67180 12788
rect 67220 12748 71788 12788
rect 71828 12748 71837 12788
rect 2563 12664 2572 12704
rect 2612 12664 2956 12704
rect 2996 12664 3005 12704
rect 4579 12664 4588 12704
rect 4628 12664 5068 12704
rect 5108 12664 5117 12704
rect 37123 12664 37132 12704
rect 37172 12664 38956 12704
rect 38996 12664 39532 12704
rect 39572 12664 39581 12704
rect 39628 12664 44812 12704
rect 44852 12664 44861 12704
rect 47875 12664 47884 12704
rect 47924 12664 48556 12704
rect 48596 12664 48605 12704
rect 48739 12664 48748 12704
rect 48788 12664 49228 12704
rect 49268 12664 49277 12704
rect 49699 12664 49708 12704
rect 49748 12664 51820 12704
rect 51860 12664 51869 12704
rect 2083 12620 2141 12621
rect 39628 12620 39668 12664
rect 53260 12620 53300 12748
rect 57283 12664 57292 12704
rect 57332 12664 58252 12704
rect 58292 12664 58301 12704
rect 62083 12664 62092 12704
rect 62132 12664 64204 12704
rect 64244 12664 64253 12704
rect 70627 12664 70636 12704
rect 70676 12664 72844 12704
rect 72884 12664 73324 12704
rect 73364 12664 73373 12704
rect 74467 12664 74476 12704
rect 74516 12664 76108 12704
rect 76148 12664 76780 12704
rect 76820 12664 76829 12704
rect 1998 12580 2092 12620
rect 2132 12580 2141 12620
rect 34915 12580 34924 12620
rect 34964 12580 39668 12620
rect 41443 12580 41452 12620
rect 41492 12580 53300 12620
rect 59299 12580 59308 12620
rect 59348 12580 61708 12620
rect 61748 12580 66892 12620
rect 66932 12580 66941 12620
rect 73987 12580 73996 12620
rect 74036 12580 74764 12620
rect 74804 12580 75820 12620
rect 75860 12580 75869 12620
rect 2083 12579 2141 12580
rect 4771 12536 4829 12537
rect 63523 12536 63581 12537
rect 63907 12536 63965 12537
rect 4483 12496 4492 12536
rect 4532 12496 4780 12536
rect 4820 12496 4829 12536
rect 36067 12496 36076 12536
rect 36116 12496 36268 12536
rect 36308 12496 36748 12536
rect 36788 12496 36797 12536
rect 38179 12496 38188 12536
rect 38228 12496 40300 12536
rect 40340 12496 40349 12536
rect 41731 12496 41740 12536
rect 41780 12496 42412 12536
rect 42452 12496 42461 12536
rect 49315 12496 49324 12536
rect 49364 12496 49612 12536
rect 49652 12496 49661 12536
rect 50947 12496 50956 12536
rect 50996 12496 51820 12536
rect 51860 12496 54412 12536
rect 54452 12496 55468 12536
rect 55508 12496 55517 12536
rect 56131 12496 56140 12536
rect 56180 12496 57580 12536
rect 57620 12496 57629 12536
rect 59011 12496 59020 12536
rect 59060 12496 59692 12536
rect 59732 12496 59741 12536
rect 63331 12496 63340 12536
rect 63380 12496 63532 12536
rect 63572 12496 63581 12536
rect 4771 12495 4829 12496
rect 63523 12495 63581 12496
rect 63628 12496 63916 12536
rect 63956 12496 64396 12536
rect 64436 12496 65548 12536
rect 65588 12496 65597 12536
rect 66019 12496 66028 12536
rect 66068 12496 68620 12536
rect 68660 12496 68669 12536
rect 69091 12496 69100 12536
rect 69140 12496 70060 12536
rect 70100 12496 70109 12536
rect 70243 12496 70252 12536
rect 70292 12496 70301 12536
rect 76387 12496 76396 12536
rect 76436 12496 76876 12536
rect 76916 12496 76925 12536
rect 77635 12496 77644 12536
rect 77684 12496 78124 12536
rect 78164 12496 78173 12536
rect 36355 12452 36413 12453
rect 63628 12452 63668 12496
rect 63907 12495 63965 12496
rect 1315 12412 1324 12452
rect 1364 12412 2996 12452
rect 36270 12412 36364 12452
rect 36404 12412 36413 12452
rect 46819 12412 46828 12452
rect 46868 12412 47020 12452
rect 47060 12412 47069 12452
rect 62275 12412 62284 12452
rect 62324 12412 63668 12452
rect 63715 12412 63724 12452
rect 63764 12412 64588 12452
rect 64628 12412 67180 12452
rect 67220 12412 67229 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 1603 12328 1612 12368
rect 1652 12328 2284 12368
rect 2324 12328 2333 12368
rect 2467 12328 2476 12368
rect 2516 12328 2860 12368
rect 2900 12328 2909 12368
rect 0 12308 80 12328
rect 1507 12244 1516 12284
rect 1556 12244 1565 12284
rect 1891 12244 1900 12284
rect 1940 12244 2188 12284
rect 2228 12244 2237 12284
rect 1516 12200 1556 12244
rect 1987 12200 2045 12201
rect 1315 12160 1324 12200
rect 1364 12160 1556 12200
rect 1699 12160 1708 12200
rect 1748 12160 1996 12200
rect 2036 12160 2045 12200
rect 1987 12159 2045 12160
rect 2956 12032 2996 12412
rect 36355 12411 36413 12412
rect 51523 12368 51581 12369
rect 5347 12328 5356 12368
rect 5396 12328 5932 12368
rect 5972 12328 5981 12368
rect 7459 12328 7468 12368
rect 7508 12328 51532 12368
rect 51572 12328 51581 12368
rect 61603 12328 61612 12368
rect 61652 12328 62092 12368
rect 62132 12328 62141 12368
rect 63235 12328 63244 12368
rect 63284 12328 64012 12368
rect 64052 12328 64340 12368
rect 51523 12327 51581 12328
rect 41827 12244 41836 12284
rect 41876 12244 42316 12284
rect 42356 12244 42365 12284
rect 45571 12244 45580 12284
rect 45620 12244 49612 12284
rect 49652 12244 49661 12284
rect 58051 12244 58060 12284
rect 58100 12244 58252 12284
rect 58292 12244 58301 12284
rect 59107 12244 59116 12284
rect 59156 12244 59404 12284
rect 59444 12244 59453 12284
rect 63043 12244 63052 12284
rect 63092 12244 63628 12284
rect 63668 12244 63677 12284
rect 36643 12200 36701 12201
rect 35011 12160 35020 12200
rect 35060 12160 36652 12200
rect 36692 12160 36701 12200
rect 36643 12159 36701 12160
rect 43180 12160 44716 12200
rect 44756 12160 53300 12200
rect 56227 12160 56236 12200
rect 56276 12160 62764 12200
rect 62804 12160 62813 12200
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 15103 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 15489 12116
rect 27103 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 27489 12116
rect 39103 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 39489 12116
rect 43180 12032 43220 12160
rect 53260 12116 53300 12160
rect 64300 12116 64340 12328
rect 70252 12200 70292 12496
rect 74563 12328 74572 12368
rect 74612 12328 74764 12368
rect 74804 12328 74813 12368
rect 78307 12244 78316 12284
rect 78356 12244 79276 12284
rect 79316 12244 79325 12284
rect 70243 12160 70252 12200
rect 70292 12160 70301 12200
rect 51103 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 51489 12116
rect 51811 12076 51820 12116
rect 51860 12076 52012 12116
rect 52052 12076 52061 12116
rect 53260 12076 59020 12116
rect 59060 12076 59069 12116
rect 63103 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 63489 12116
rect 64300 12076 64396 12116
rect 64436 12076 64445 12116
rect 69667 12076 69676 12116
rect 69716 12076 70348 12116
rect 70388 12076 70397 12116
rect 75103 12076 75112 12116
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75480 12076 75489 12116
rect 2956 11992 3476 12032
rect 42403 11992 42412 12032
rect 42452 11992 43220 12032
rect 44611 11992 44620 12032
rect 44660 11992 46828 12032
rect 46868 11992 46877 12032
rect 57475 11992 57484 12032
rect 57524 11992 66220 12032
rect 66260 11992 66269 12032
rect 69955 11992 69964 12032
rect 70004 11992 70540 12032
rect 70580 11992 70589 12032
rect 3436 11948 3476 11992
rect 52195 11948 52253 11949
rect 57484 11948 57524 11992
rect 3427 11908 3436 11948
rect 3476 11908 3485 11948
rect 33859 11908 33868 11948
rect 33908 11908 34828 11948
rect 34868 11908 34877 11948
rect 45475 11908 45484 11948
rect 45524 11908 48268 11948
rect 48308 11908 48317 11948
rect 50275 11908 50284 11948
rect 50324 11908 50764 11948
rect 50804 11908 50813 11948
rect 52195 11908 52204 11948
rect 52244 11908 57524 11948
rect 60643 11948 60701 11949
rect 60643 11908 60652 11948
rect 60692 11908 61036 11948
rect 61076 11908 61085 11948
rect 62563 11908 62572 11948
rect 62612 11908 62764 11948
rect 62804 11908 63244 11948
rect 63284 11908 63532 11948
rect 63572 11908 63581 11948
rect 69475 11908 69484 11948
rect 69524 11908 69868 11948
rect 69908 11908 69917 11948
rect 74947 11908 74956 11948
rect 74996 11908 75724 11948
rect 75764 11908 75773 11948
rect 2083 11864 2141 11865
rect 50764 11864 50804 11908
rect 52195 11907 52253 11908
rect 60643 11907 60701 11908
rect 1998 11824 2092 11864
rect 2132 11824 2141 11864
rect 3331 11824 3340 11864
rect 3380 11824 3532 11864
rect 3572 11824 3916 11864
rect 3956 11824 3965 11864
rect 44515 11824 44524 11864
rect 44564 11824 44908 11864
rect 44948 11824 44957 11864
rect 48547 11824 48556 11864
rect 48596 11824 49132 11864
rect 49172 11824 49181 11864
rect 50764 11824 52204 11864
rect 52244 11824 52253 11864
rect 60739 11824 60748 11864
rect 60788 11824 63380 11864
rect 63427 11824 63436 11864
rect 63476 11824 64204 11864
rect 64244 11824 64876 11864
rect 64916 11824 64925 11864
rect 68803 11824 68812 11864
rect 68852 11824 69004 11864
rect 69044 11824 70060 11864
rect 70100 11824 73460 11864
rect 2083 11823 2141 11824
rect 47683 11780 47741 11781
rect 63340 11780 63380 11824
rect 73420 11780 73460 11824
rect 1411 11740 1420 11780
rect 1460 11740 7468 11780
rect 7508 11740 7517 11780
rect 38860 11740 41452 11780
rect 41492 11740 41501 11780
rect 46531 11740 46540 11780
rect 46580 11740 47692 11780
rect 47732 11740 47741 11780
rect 50371 11740 50380 11780
rect 50420 11740 51860 11780
rect 56803 11740 56812 11780
rect 56852 11740 57964 11780
rect 58004 11740 58156 11780
rect 58196 11740 58205 11780
rect 58339 11740 58348 11780
rect 58388 11740 62572 11780
rect 62612 11740 62621 11780
rect 63340 11740 64588 11780
rect 64628 11740 64972 11780
rect 65012 11740 65452 11780
rect 65492 11740 65501 11780
rect 69859 11740 69868 11780
rect 69908 11740 70636 11780
rect 70676 11740 70685 11780
rect 73420 11740 73996 11780
rect 74036 11740 74045 11780
rect 75628 11740 77068 11780
rect 77108 11740 78316 11780
rect 78356 11740 78365 11780
rect 38860 11696 38900 11740
rect 47683 11739 47741 11740
rect 1987 11656 1996 11696
rect 2036 11656 2668 11696
rect 2708 11656 3724 11696
rect 3764 11656 3916 11696
rect 3956 11656 3965 11696
rect 34819 11656 34828 11696
rect 34868 11656 35308 11696
rect 35348 11656 35357 11696
rect 35587 11656 35596 11696
rect 35636 11656 36076 11696
rect 36116 11656 36125 11696
rect 38851 11656 38860 11696
rect 38900 11656 38909 11696
rect 39139 11656 39148 11696
rect 39188 11656 39532 11696
rect 39572 11656 39581 11696
rect 43555 11656 43564 11696
rect 43604 11656 44332 11696
rect 44372 11656 45388 11696
rect 45428 11656 45437 11696
rect 46915 11656 46924 11696
rect 46964 11656 47116 11696
rect 47156 11656 47165 11696
rect 48451 11656 48460 11696
rect 48500 11656 49228 11696
rect 49268 11656 49277 11696
rect 49411 11656 49420 11696
rect 49460 11656 50228 11696
rect 50188 11612 50228 11656
rect 51820 11612 51860 11740
rect 68899 11696 68957 11697
rect 75628 11696 75668 11740
rect 51907 11656 51916 11696
rect 51956 11656 52108 11696
rect 52148 11656 53356 11696
rect 53396 11656 53405 11696
rect 53923 11656 53932 11696
rect 53972 11656 56236 11696
rect 56276 11656 56285 11696
rect 58819 11656 58828 11696
rect 58868 11656 60748 11696
rect 60788 11656 60797 11696
rect 62083 11656 62092 11696
rect 62132 11656 66028 11696
rect 66068 11656 66077 11696
rect 68814 11656 68908 11696
rect 68948 11656 68957 11696
rect 69283 11656 69292 11696
rect 69332 11656 70444 11696
rect 70484 11656 70493 11696
rect 75619 11656 75628 11696
rect 75668 11656 75677 11696
rect 76195 11656 76204 11696
rect 76244 11656 76588 11696
rect 76628 11656 76637 11696
rect 68899 11655 68957 11656
rect 70531 11612 70589 11613
rect 76204 11612 76244 11656
rect 3619 11572 3628 11612
rect 3668 11572 5068 11612
rect 5108 11572 7372 11612
rect 7412 11572 34924 11612
rect 34964 11572 34973 11612
rect 36835 11572 36844 11612
rect 36884 11572 37996 11612
rect 38036 11572 39340 11612
rect 39380 11572 39389 11612
rect 50179 11572 50188 11612
rect 50228 11572 51148 11612
rect 51188 11572 51197 11612
rect 51820 11572 52148 11612
rect 57283 11572 57292 11612
rect 57332 11572 58348 11612
rect 58388 11572 58397 11612
rect 58915 11572 58924 11612
rect 58964 11572 59308 11612
rect 59348 11572 59357 11612
rect 62755 11572 62764 11612
rect 62804 11572 63820 11612
rect 63860 11572 63869 11612
rect 67363 11572 67372 11612
rect 67412 11572 69004 11612
rect 69044 11572 69053 11612
rect 70243 11572 70252 11612
rect 70292 11572 70540 11612
rect 70580 11572 70589 11612
rect 0 11528 80 11548
rect 50380 11528 50420 11572
rect 52108 11528 52148 11572
rect 70531 11571 70589 11572
rect 75340 11572 76244 11612
rect 76387 11612 76445 11613
rect 76387 11572 76396 11612
rect 76436 11572 77164 11612
rect 77204 11572 77213 11612
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 4195 11488 4204 11528
rect 4244 11488 4684 11528
rect 4724 11488 4733 11528
rect 36451 11488 36460 11528
rect 36500 11488 38188 11528
rect 38228 11488 39628 11528
rect 39668 11488 39677 11528
rect 49123 11488 49132 11528
rect 49172 11488 49804 11528
rect 49844 11488 49853 11528
rect 50371 11488 50380 11528
rect 50420 11488 50429 11528
rect 52099 11488 52108 11528
rect 52148 11488 52157 11528
rect 59491 11488 59500 11528
rect 59540 11488 60844 11528
rect 60884 11488 63764 11528
rect 0 11468 80 11488
rect 63724 11444 63764 11488
rect 3427 11404 3436 11444
rect 3476 11404 3628 11444
rect 3668 11404 3677 11444
rect 35491 11404 35500 11444
rect 35540 11404 37036 11444
rect 37076 11404 37085 11444
rect 61795 11404 61804 11444
rect 61844 11404 63436 11444
rect 63476 11404 63485 11444
rect 63724 11404 63916 11444
rect 63956 11404 63965 11444
rect 74851 11360 74909 11361
rect 75340 11360 75380 11572
rect 76387 11571 76445 11572
rect 75427 11488 75436 11528
rect 75476 11488 76012 11528
rect 76052 11488 76061 11528
rect 76204 11488 76300 11528
rect 76340 11488 76349 11528
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 16343 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 16729 11360
rect 28343 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 28729 11360
rect 40343 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 40729 11360
rect 42115 11320 42124 11360
rect 42164 11320 43220 11360
rect 52343 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 52729 11360
rect 63235 11320 63244 11360
rect 63284 11320 63820 11360
rect 63860 11320 63869 11360
rect 64343 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 64729 11360
rect 74766 11320 74860 11360
rect 74900 11320 74909 11360
rect 75331 11320 75340 11360
rect 75380 11320 75389 11360
rect 43180 11276 43220 11320
rect 74851 11319 74909 11320
rect 76204 11276 76244 11488
rect 76343 11320 76352 11360
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76720 11320 76729 11360
rect 43180 11236 43948 11276
rect 43988 11236 46252 11276
rect 46292 11236 46301 11276
rect 70339 11236 70348 11276
rect 70388 11236 76340 11276
rect 4771 11192 4829 11193
rect 76300 11192 76340 11236
rect 4579 11152 4588 11192
rect 4628 11152 4780 11192
rect 4820 11152 4829 11192
rect 42115 11152 42124 11192
rect 42164 11152 42508 11192
rect 42548 11152 42557 11192
rect 43459 11152 43468 11192
rect 43508 11152 43852 11192
rect 43892 11152 46540 11192
rect 46580 11152 46589 11192
rect 58435 11152 58444 11192
rect 58484 11152 58828 11192
rect 58868 11152 59308 11192
rect 59348 11152 59357 11192
rect 60931 11152 60940 11192
rect 60980 11152 62380 11192
rect 62420 11152 62764 11192
rect 62804 11152 62813 11192
rect 72451 11152 72460 11192
rect 72500 11152 75244 11192
rect 75284 11152 75293 11192
rect 76291 11152 76300 11192
rect 76340 11152 77260 11192
rect 77300 11152 77309 11192
rect 4771 11151 4829 11152
rect 3811 11068 3820 11108
rect 3860 11068 4300 11108
rect 4340 11068 4349 11108
rect 48067 11068 48076 11108
rect 48116 11068 50860 11108
rect 50900 11068 50909 11108
rect 53260 11068 53740 11108
rect 53780 11068 53789 11108
rect 69667 11068 69676 11108
rect 69716 11068 70156 11108
rect 70196 11068 70205 11108
rect 4867 11024 4925 11025
rect 40867 11024 40925 11025
rect 49315 11024 49373 11025
rect 53260 11024 53300 11068
rect 4782 10984 4876 11024
rect 4916 10984 4925 11024
rect 35395 10984 35404 11024
rect 35444 10984 36940 11024
rect 36980 10984 36989 11024
rect 37123 10984 37132 11024
rect 37172 10984 38764 11024
rect 38804 10984 38813 11024
rect 39427 10984 39436 11024
rect 39476 10984 40876 11024
rect 40916 10984 44564 11024
rect 49230 10984 49324 11024
rect 49364 10984 49373 11024
rect 49987 10984 49996 11024
rect 50036 10984 51340 11024
rect 51380 10984 53300 11024
rect 53347 10984 53356 11024
rect 53396 10984 54124 11024
rect 54164 10984 54173 11024
rect 59683 10984 59692 11024
rect 59732 10984 61804 11024
rect 61844 10984 61853 11024
rect 62179 10984 62188 11024
rect 62228 10984 62956 11024
rect 62996 10984 63005 11024
rect 63907 10984 63916 11024
rect 63956 10984 64588 11024
rect 64628 10984 64637 11024
rect 74659 10984 74668 11024
rect 74708 10984 75148 11024
rect 75188 10984 75197 11024
rect 75811 10984 75820 11024
rect 75860 10984 76684 11024
rect 76724 10984 76733 11024
rect 4867 10983 4925 10984
rect 40867 10983 40925 10984
rect 36163 10816 36172 10856
rect 36212 10816 36748 10856
rect 36788 10816 36797 10856
rect 41539 10816 41548 10856
rect 41588 10816 43084 10856
rect 43124 10816 43133 10856
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 40003 10732 40012 10772
rect 40052 10732 42028 10772
rect 42068 10732 42508 10772
rect 42548 10732 42557 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 44524 10688 44564 10984
rect 49315 10983 49373 10984
rect 64675 10900 64684 10940
rect 64724 10900 65164 10940
rect 65204 10900 65213 10940
rect 46531 10816 46540 10856
rect 46580 10816 60076 10856
rect 60116 10816 60125 10856
rect 53347 10732 53356 10772
rect 53396 10732 53836 10772
rect 53876 10732 53885 10772
rect 70723 10732 70732 10772
rect 70772 10732 71116 10772
rect 71156 10732 71165 10772
rect 44524 10648 50668 10688
rect 50708 10648 50717 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 15103 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 15489 10604
rect 27103 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 27489 10604
rect 38851 10564 38860 10604
rect 38900 10564 38909 10604
rect 39103 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 39489 10604
rect 51103 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 51489 10604
rect 63103 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 63489 10604
rect 68899 10564 68908 10604
rect 68948 10564 69388 10604
rect 69428 10564 69437 10604
rect 75103 10564 75112 10604
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75480 10564 75489 10604
rect 1315 10396 1324 10436
rect 1364 10396 3436 10436
rect 3476 10396 3485 10436
rect 38860 10352 38900 10564
rect 53260 10480 60364 10520
rect 60404 10480 60413 10520
rect 68419 10480 68428 10520
rect 68468 10480 69484 10520
rect 69524 10480 69533 10520
rect 53260 10436 53300 10480
rect 63523 10436 63581 10437
rect 42115 10396 42124 10436
rect 42164 10396 43220 10436
rect 46819 10396 46828 10436
rect 46868 10396 47116 10436
rect 47156 10396 49132 10436
rect 49172 10396 53300 10436
rect 56419 10396 56428 10436
rect 56468 10396 58060 10436
rect 58100 10396 58109 10436
rect 63427 10396 63436 10436
rect 63476 10396 63532 10436
rect 63572 10396 63581 10436
rect 64579 10396 64588 10436
rect 64628 10396 65452 10436
rect 65492 10396 67660 10436
rect 67700 10396 71500 10436
rect 71540 10396 71549 10436
rect 72835 10396 72844 10436
rect 72884 10396 73516 10436
rect 73556 10396 73565 10436
rect 75907 10396 75916 10436
rect 75956 10396 76588 10436
rect 76628 10396 76637 10436
rect 43180 10352 43220 10396
rect 63523 10395 63581 10396
rect 931 10312 940 10352
rect 980 10312 1516 10352
rect 1556 10312 1565 10352
rect 1612 10312 2188 10352
rect 2228 10312 2237 10352
rect 2467 10312 2476 10352
rect 2516 10312 2668 10352
rect 2708 10312 2717 10352
rect 5059 10312 5068 10352
rect 5108 10312 5260 10352
rect 5300 10312 5309 10352
rect 38860 10312 39188 10352
rect 43180 10312 48364 10352
rect 48404 10312 48413 10352
rect 50275 10312 50284 10352
rect 50324 10312 52012 10352
rect 52052 10312 52061 10352
rect 57571 10312 57580 10352
rect 57620 10312 58252 10352
rect 58292 10312 58301 10352
rect 58732 10312 61996 10352
rect 62036 10312 63476 10352
rect 67267 10312 67276 10352
rect 67316 10312 67852 10352
rect 67892 10312 67901 10352
rect 68899 10312 68908 10352
rect 68948 10312 69772 10352
rect 69812 10312 70060 10352
rect 70100 10312 70109 10352
rect 1612 10268 1652 10312
rect 39148 10268 39188 10312
rect 58732 10268 58772 10312
rect 58915 10268 58973 10269
rect 1603 10228 1612 10268
rect 1652 10228 1661 10268
rect 3331 10228 3340 10268
rect 3380 10228 4876 10268
rect 4916 10228 4925 10268
rect 39139 10228 39148 10268
rect 39188 10228 39197 10268
rect 46243 10228 46252 10268
rect 46292 10228 48844 10268
rect 48884 10228 48893 10268
rect 57379 10228 57388 10268
rect 57428 10228 58732 10268
rect 58772 10228 58781 10268
rect 58830 10228 58924 10268
rect 58964 10228 58973 10268
rect 58915 10227 58973 10228
rect 63436 10184 63476 10312
rect 68227 10228 68236 10268
rect 68276 10228 68620 10268
rect 68660 10228 68669 10268
rect 69283 10228 69292 10268
rect 69332 10228 70636 10268
rect 70676 10228 70685 10268
rect 76483 10228 76492 10268
rect 76532 10228 77740 10268
rect 77780 10228 79468 10268
rect 79508 10228 79517 10268
rect 2371 10144 2380 10184
rect 2420 10144 4204 10184
rect 4244 10144 4253 10184
rect 43075 10144 43084 10184
rect 43124 10144 43468 10184
rect 43508 10144 46964 10184
rect 52963 10144 52972 10184
rect 53012 10144 53932 10184
rect 53972 10144 53981 10184
rect 57859 10144 57868 10184
rect 57908 10144 59212 10184
rect 59252 10144 59261 10184
rect 59884 10144 63380 10184
rect 63427 10144 63436 10184
rect 63476 10144 64204 10184
rect 64244 10144 64253 10184
rect 68515 10144 68524 10184
rect 68564 10144 69196 10184
rect 69236 10144 69676 10184
rect 69716 10144 69725 10184
rect 70819 10144 70828 10184
rect 70868 10144 71308 10184
rect 71348 10144 71357 10184
rect 71683 10144 71692 10184
rect 71732 10144 72940 10184
rect 72980 10144 74668 10184
rect 74708 10144 78316 10184
rect 78356 10144 78365 10184
rect 2851 10060 2860 10100
rect 2900 10060 3148 10100
rect 3188 10060 3197 10100
rect 38659 10060 38668 10100
rect 38708 10060 39244 10100
rect 39284 10060 39293 10100
rect 40867 10060 40876 10100
rect 40916 10060 41740 10100
rect 41780 10060 41789 10100
rect 42211 10060 42220 10100
rect 42260 10060 43660 10100
rect 43700 10060 44428 10100
rect 44468 10060 44477 10100
rect 46339 10060 46348 10100
rect 46388 10060 46732 10100
rect 46772 10060 46781 10100
rect 4771 10016 4829 10017
rect 4579 9976 4588 10016
rect 4628 9976 4780 10016
rect 4820 9976 4829 10016
rect 40579 9976 40588 10016
rect 40628 9976 41836 10016
rect 41876 9976 41885 10016
rect 4771 9975 4829 9976
rect 46924 9932 46964 10144
rect 59884 10100 59924 10144
rect 63340 10100 63380 10144
rect 69091 10100 69149 10101
rect 53155 10060 53164 10100
rect 53204 10060 53644 10100
rect 53684 10060 53693 10100
rect 59875 10060 59884 10100
rect 59924 10060 59933 10100
rect 63340 10060 63628 10100
rect 63668 10060 65164 10100
rect 65204 10060 65213 10100
rect 66883 10060 66892 10100
rect 66932 10060 68812 10100
rect 68852 10060 68861 10100
rect 69006 10060 69100 10100
rect 69140 10060 69149 10100
rect 69571 10060 69580 10100
rect 69620 10060 72844 10100
rect 72884 10060 72893 10100
rect 73411 10060 73420 10100
rect 73460 10060 75916 10100
rect 75956 10060 75965 10100
rect 76291 10060 76300 10100
rect 76340 10060 76876 10100
rect 76916 10060 76925 10100
rect 69091 10059 69149 10060
rect 70924 10016 70964 10060
rect 52291 9976 52300 10016
rect 52340 9976 52349 10016
rect 52675 9976 52684 10016
rect 52724 9976 53452 10016
rect 53492 9976 53501 10016
rect 58051 9976 58060 10016
rect 58100 9976 58348 10016
rect 58388 9976 58397 10016
rect 59971 9976 59980 10016
rect 60020 9976 60268 10016
rect 60308 9976 60317 10016
rect 70915 9976 70924 10016
rect 70964 9976 70973 10016
rect 76204 9976 76396 10016
rect 76436 9976 76445 10016
rect 52300 9932 52340 9976
rect 41740 9892 42316 9932
rect 42356 9892 43276 9932
rect 43316 9892 43325 9932
rect 46915 9892 46924 9932
rect 46964 9892 46973 9932
rect 52300 9892 53068 9932
rect 53108 9892 53117 9932
rect 68323 9892 68332 9932
rect 68372 9892 69676 9932
rect 69716 9892 69725 9932
rect 71107 9892 71116 9932
rect 71156 9892 71692 9932
rect 71732 9892 71741 9932
rect 0 9848 80 9868
rect 41740 9848 41780 9892
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 16343 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 16729 9848
rect 28343 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 28729 9848
rect 40343 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 40729 9848
rect 41731 9808 41740 9848
rect 41780 9808 41789 9848
rect 52343 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 52729 9848
rect 64343 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 64729 9848
rect 75523 9808 75532 9848
rect 75572 9808 76012 9848
rect 76052 9808 76061 9848
rect 0 9788 80 9808
rect 48643 9764 48701 9765
rect 76204 9764 76244 9976
rect 76343 9808 76352 9848
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76720 9808 76729 9848
rect 7171 9724 7180 9764
rect 7220 9724 48652 9764
rect 48692 9724 48701 9764
rect 72547 9724 72556 9764
rect 72596 9724 76532 9764
rect 48643 9723 48701 9724
rect 76492 9680 76532 9724
rect 835 9640 844 9680
rect 884 9640 1516 9680
rect 1556 9640 1565 9680
rect 2851 9640 2860 9680
rect 2900 9640 3532 9680
rect 3572 9640 3581 9680
rect 39331 9640 39340 9680
rect 39380 9640 40108 9680
rect 40148 9640 40157 9680
rect 40771 9640 40780 9680
rect 40820 9640 42796 9680
rect 42836 9640 43084 9680
rect 43124 9640 43133 9680
rect 49891 9640 49900 9680
rect 49940 9640 53068 9680
rect 53108 9640 53117 9680
rect 61987 9640 61996 9680
rect 62036 9640 66796 9680
rect 66836 9640 66845 9680
rect 74851 9640 74860 9680
rect 74900 9640 75724 9680
rect 75764 9640 75773 9680
rect 76483 9640 76492 9680
rect 76532 9640 76541 9680
rect 77347 9640 77356 9680
rect 77396 9640 78124 9680
rect 78164 9640 79468 9680
rect 79508 9640 79517 9680
rect 76195 9596 76253 9597
rect 77356 9596 77396 9640
rect 3619 9556 3628 9596
rect 3668 9556 3677 9596
rect 4483 9556 4492 9596
rect 4532 9556 4780 9596
rect 4820 9556 4829 9596
rect 40675 9556 40684 9596
rect 40724 9556 41356 9596
rect 41396 9556 41405 9596
rect 41923 9556 41932 9596
rect 41972 9556 42988 9596
rect 43028 9556 43037 9596
rect 52099 9556 52108 9596
rect 52148 9556 52396 9596
rect 52436 9556 52445 9596
rect 62179 9556 62188 9596
rect 62228 9556 64876 9596
rect 64916 9556 64925 9596
rect 69859 9556 69868 9596
rect 69908 9556 71212 9596
rect 71252 9556 71261 9596
rect 74563 9556 74572 9596
rect 74612 9556 75628 9596
rect 75668 9556 76204 9596
rect 76244 9556 76253 9596
rect 76579 9556 76588 9596
rect 76628 9556 77396 9596
rect 1987 9472 1996 9512
rect 2036 9472 2956 9512
rect 2996 9472 3244 9512
rect 3284 9472 3293 9512
rect 3628 9428 3668 9556
rect 41356 9512 41396 9556
rect 4291 9472 4300 9512
rect 4340 9472 4876 9512
rect 4916 9472 4925 9512
rect 29155 9472 29164 9512
rect 29204 9472 39436 9512
rect 39476 9472 39485 9512
rect 40195 9472 40204 9512
rect 40244 9472 40588 9512
rect 40628 9472 40637 9512
rect 41356 9472 42700 9512
rect 42740 9472 42749 9512
rect 42883 9472 42892 9512
rect 42932 9472 43852 9512
rect 43892 9472 43901 9512
rect 44515 9472 44524 9512
rect 44564 9472 45868 9512
rect 45908 9472 48460 9512
rect 48500 9472 48509 9512
rect 53731 9472 53740 9512
rect 53780 9472 54508 9512
rect 54548 9472 54557 9512
rect 60835 9472 60844 9512
rect 60884 9472 63436 9512
rect 63476 9472 66604 9512
rect 66644 9472 66653 9512
rect 70147 9472 70156 9512
rect 70196 9472 70828 9512
rect 70868 9472 70877 9512
rect 71107 9472 71116 9512
rect 71156 9472 71884 9512
rect 71924 9472 74092 9512
rect 74132 9472 74141 9512
rect 42700 9428 42740 9472
rect 835 9388 844 9428
rect 884 9388 1420 9428
rect 1460 9388 1469 9428
rect 3139 9388 3148 9428
rect 3188 9388 4492 9428
rect 4532 9388 4541 9428
rect 42700 9388 45388 9428
rect 45428 9388 45437 9428
rect 69379 9388 69388 9428
rect 69428 9388 70580 9428
rect 71683 9388 71692 9428
rect 71732 9388 72556 9428
rect 72596 9388 72605 9428
rect 4771 9344 4829 9345
rect 70540 9344 70580 9388
rect 74764 9344 74804 9556
rect 76195 9555 76253 9556
rect 76195 9472 76204 9512
rect 76244 9472 77260 9512
rect 77300 9472 77309 9512
rect 77356 9472 77548 9512
rect 77588 9472 77932 9512
rect 77972 9472 77981 9512
rect 77356 9428 77396 9472
rect 76771 9388 76780 9428
rect 76820 9388 77396 9428
rect 4579 9304 4588 9344
rect 4628 9304 4780 9344
rect 4820 9304 4829 9344
rect 43075 9304 43084 9344
rect 43124 9304 45580 9344
rect 45620 9304 45629 9344
rect 58627 9304 58636 9344
rect 58676 9304 60212 9344
rect 69859 9304 69868 9344
rect 69908 9304 70444 9344
rect 70484 9304 70493 9344
rect 70540 9304 74804 9344
rect 4771 9303 4829 9304
rect 60172 9260 60212 9304
rect 3427 9220 3436 9260
rect 3476 9220 3628 9260
rect 3668 9220 3677 9260
rect 41539 9220 41548 9260
rect 41588 9220 42412 9260
rect 42452 9220 42461 9260
rect 44899 9220 44908 9260
rect 44948 9220 45964 9260
rect 46004 9220 46444 9260
rect 46484 9220 46493 9260
rect 52675 9220 52684 9260
rect 52724 9220 59308 9260
rect 59348 9220 59357 9260
rect 60163 9220 60172 9260
rect 60212 9220 61996 9260
rect 62036 9220 62045 9260
rect 63811 9220 63820 9260
rect 63860 9220 64588 9260
rect 64628 9220 64637 9260
rect 68899 9220 68908 9260
rect 68948 9220 71404 9260
rect 71444 9220 71884 9260
rect 71924 9220 71933 9260
rect 75811 9220 75820 9260
rect 75860 9220 76684 9260
rect 76724 9220 76733 9260
rect 77356 9176 77396 9388
rect 49891 9136 49900 9176
rect 49940 9136 50764 9176
rect 50804 9136 57196 9176
rect 57236 9136 57245 9176
rect 58339 9136 58348 9176
rect 58388 9136 59212 9176
rect 59252 9136 60364 9176
rect 60404 9136 60413 9176
rect 70540 9136 71308 9176
rect 71348 9136 71357 9176
rect 77347 9136 77356 9176
rect 77396 9136 77405 9176
rect 70540 9092 70580 9136
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 15103 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 15489 9092
rect 27103 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 27489 9092
rect 39103 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 39489 9092
rect 51103 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 51489 9092
rect 58051 9052 58060 9092
rect 58100 9052 58252 9092
rect 58292 9052 58732 9092
rect 58772 9052 58781 9092
rect 59299 9052 59308 9092
rect 59348 9052 59884 9092
rect 59924 9052 59933 9092
rect 63103 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 63489 9092
rect 70531 9052 70540 9092
rect 70580 9052 70589 9092
rect 75103 9052 75112 9092
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75480 9052 75489 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 53260 8968 53452 9008
rect 53492 8968 53501 9008
rect 53548 8968 54220 9008
rect 54260 8968 56812 9008
rect 56852 8968 62668 9008
rect 62708 8968 62717 9008
rect 64099 8968 64108 9008
rect 64148 8968 64780 9008
rect 64820 8968 64829 9008
rect 69283 8968 69292 9008
rect 69332 8968 69676 9008
rect 69716 8968 69725 9008
rect 0 8948 80 8968
rect 53260 8924 53300 8968
rect 53548 8924 53588 8968
rect 51340 8884 51916 8924
rect 51956 8884 52684 8924
rect 52724 8884 52733 8924
rect 53251 8884 53260 8924
rect 53300 8884 53309 8924
rect 53539 8884 53548 8924
rect 53588 8884 53597 8924
rect 59011 8884 59020 8924
rect 59060 8884 59692 8924
rect 59732 8884 59741 8924
rect 2755 8800 2764 8840
rect 2804 8800 3436 8840
rect 3476 8800 3485 8840
rect 4771 8800 4780 8840
rect 4820 8800 4972 8840
rect 5012 8800 5021 8840
rect 47980 8800 49228 8840
rect 49268 8800 49277 8840
rect 47980 8756 48020 8800
rect 1228 8716 1996 8756
rect 2036 8716 3532 8756
rect 3572 8716 3581 8756
rect 41827 8716 41836 8756
rect 41876 8716 42796 8756
rect 42836 8716 45484 8756
rect 45524 8716 46540 8756
rect 46580 8716 47980 8756
rect 48020 8716 48029 8756
rect 48163 8716 48172 8756
rect 48212 8716 48460 8756
rect 48500 8716 48509 8756
rect 1228 8588 1268 8716
rect 51340 8672 51380 8884
rect 51523 8800 51532 8840
rect 51572 8800 51820 8840
rect 51860 8800 52876 8840
rect 52916 8800 53740 8840
rect 53780 8800 54028 8840
rect 54068 8800 54412 8840
rect 54452 8800 54461 8840
rect 57763 8800 57772 8840
rect 57812 8800 57821 8840
rect 57955 8800 57964 8840
rect 58004 8800 58013 8840
rect 58252 8800 58540 8840
rect 58580 8800 62860 8840
rect 62900 8800 62909 8840
rect 64387 8800 64396 8840
rect 64436 8800 65068 8840
rect 65108 8800 65117 8840
rect 68995 8800 69004 8840
rect 69044 8800 69196 8840
rect 69236 8800 69245 8840
rect 69379 8800 69388 8840
rect 69428 8800 70156 8840
rect 70196 8800 70732 8840
rect 70772 8800 70781 8840
rect 51619 8716 51628 8756
rect 51668 8716 52204 8756
rect 52244 8716 52253 8756
rect 1699 8632 1708 8672
rect 1748 8632 2900 8672
rect 4483 8632 4492 8672
rect 4532 8632 4972 8672
rect 5012 8632 7180 8672
rect 7220 8632 7229 8672
rect 41443 8632 41452 8672
rect 41492 8632 41932 8672
rect 41972 8632 41981 8672
rect 49123 8632 49132 8672
rect 49172 8632 49804 8672
rect 49844 8632 49853 8672
rect 49987 8632 49996 8672
rect 50036 8632 51340 8672
rect 51380 8632 51389 8672
rect 51820 8632 52108 8672
rect 52148 8632 52157 8672
rect 52387 8632 52396 8672
rect 52436 8632 53164 8672
rect 53204 8632 53213 8672
rect 53443 8632 53452 8672
rect 53492 8632 53932 8672
rect 53972 8632 53981 8672
rect 2860 8588 2900 8632
rect 51820 8588 51860 8632
rect 57772 8588 57812 8800
rect 57964 8672 58004 8800
rect 58252 8756 58292 8800
rect 58243 8716 58252 8756
rect 58292 8716 58301 8756
rect 59308 8716 59692 8756
rect 59732 8716 59741 8756
rect 59308 8672 59348 8716
rect 57964 8632 59348 8672
rect 59395 8632 59404 8672
rect 59444 8632 60076 8672
rect 60116 8632 60125 8672
rect 62851 8632 62860 8672
rect 62900 8632 64012 8672
rect 64052 8632 64061 8672
rect 66595 8632 66604 8672
rect 66644 8632 67276 8672
rect 67316 8632 68140 8672
rect 68180 8632 68189 8672
rect 68707 8632 68716 8672
rect 68756 8632 69580 8672
rect 69620 8632 69629 8672
rect 59308 8588 59348 8632
rect 1219 8548 1228 8588
rect 1268 8548 1277 8588
rect 2860 8548 7700 8588
rect 46915 8548 46924 8588
rect 46964 8548 47980 8588
rect 48020 8548 48029 8588
rect 48547 8548 48556 8588
rect 48596 8548 49036 8588
rect 49076 8548 49085 8588
rect 50179 8548 50188 8588
rect 50228 8548 51860 8588
rect 51916 8548 55084 8588
rect 55124 8548 55660 8588
rect 55700 8548 55709 8588
rect 55939 8548 55948 8588
rect 55988 8548 57812 8588
rect 59299 8548 59308 8588
rect 59348 8548 59357 8588
rect 69187 8548 69196 8588
rect 69236 8548 70060 8588
rect 70100 8548 70109 8588
rect 75715 8548 75724 8588
rect 75764 8548 76300 8588
rect 76340 8548 76349 8588
rect 76579 8548 76588 8588
rect 76628 8548 76637 8588
rect 7660 8504 7700 8548
rect 50851 8504 50909 8505
rect 51916 8504 51956 8548
rect 76588 8504 76628 8548
rect 2467 8464 2476 8504
rect 2516 8464 3820 8504
rect 3860 8464 4396 8504
rect 4436 8464 4445 8504
rect 7651 8464 7660 8504
rect 7700 8464 50860 8504
rect 50900 8464 50909 8504
rect 51715 8464 51724 8504
rect 51764 8464 51956 8504
rect 52771 8464 52780 8504
rect 52820 8464 53356 8504
rect 53396 8464 53405 8504
rect 57859 8464 57868 8504
rect 57908 8464 58444 8504
rect 58484 8464 58732 8504
rect 58772 8464 58781 8504
rect 60259 8464 60268 8504
rect 60308 8464 60317 8504
rect 64483 8464 64492 8504
rect 64532 8464 64876 8504
rect 64916 8464 64925 8504
rect 69667 8464 69676 8504
rect 69716 8464 70348 8504
rect 70388 8464 70397 8504
rect 75907 8464 75916 8504
rect 75956 8464 76628 8504
rect 50851 8463 50909 8464
rect 60268 8420 60308 8464
rect 76195 8420 76253 8421
rect 52963 8380 52972 8420
rect 53012 8380 53644 8420
rect 53684 8380 53693 8420
rect 55171 8380 55180 8420
rect 55220 8380 60308 8420
rect 76110 8380 76204 8420
rect 76244 8380 76253 8420
rect 76195 8379 76253 8380
rect 48835 8336 48893 8337
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 16343 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 16729 8336
rect 28343 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 28729 8336
rect 40343 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 40729 8336
rect 48750 8296 48844 8336
rect 48884 8296 48893 8336
rect 52343 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 52729 8336
rect 59299 8296 59308 8336
rect 59348 8296 59980 8336
rect 60020 8296 60029 8336
rect 64343 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 64729 8336
rect 68419 8296 68428 8336
rect 68468 8296 71020 8336
rect 71060 8296 71069 8336
rect 76343 8296 76352 8336
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76720 8296 76729 8336
rect 48835 8295 48893 8296
rect 48259 8212 48268 8252
rect 48308 8212 49900 8252
rect 49940 8212 49949 8252
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 1123 8128 1132 8168
rect 1172 8128 2380 8168
rect 2420 8128 2429 8168
rect 44227 8128 44236 8168
rect 44276 8128 45004 8168
rect 45044 8128 45053 8168
rect 48748 8128 48940 8168
rect 48980 8128 48989 8168
rect 60067 8128 60076 8168
rect 60116 8128 62860 8168
rect 62900 8128 67756 8168
rect 67796 8128 67805 8168
rect 75907 8128 75916 8168
rect 75956 8128 76396 8168
rect 76436 8128 76445 8168
rect 0 8108 80 8128
rect 42979 8044 42988 8084
rect 43028 8044 44468 8084
rect 4771 8000 4829 8001
rect 44428 8000 44468 8044
rect 1795 7960 1804 8000
rect 1844 7960 3052 8000
rect 3092 7960 3820 8000
rect 3860 7960 3869 8000
rect 4579 7960 4588 8000
rect 4628 7960 4780 8000
rect 4820 7960 6412 8000
rect 6452 7960 6461 8000
rect 44419 7960 44428 8000
rect 44468 7960 44477 8000
rect 45667 7960 45676 8000
rect 45716 7960 46732 8000
rect 46772 7960 46781 8000
rect 47011 7960 47020 8000
rect 47060 7960 47069 8000
rect 47299 7960 47308 8000
rect 47348 7960 48556 8000
rect 48596 7960 48605 8000
rect 4771 7959 4829 7960
rect 44428 7916 44468 7960
rect 47020 7916 47060 7960
rect 44428 7876 47692 7916
rect 47732 7876 47741 7916
rect 48748 7832 48788 8128
rect 52195 8044 52204 8084
rect 52244 8044 52684 8084
rect 52724 8044 53260 8084
rect 53300 8044 53309 8084
rect 74851 8044 74860 8084
rect 74900 8044 76300 8084
rect 76340 8044 76349 8084
rect 66307 8000 66365 8001
rect 48835 7960 48844 8000
rect 48884 7960 49228 8000
rect 49268 7960 49277 8000
rect 53260 7960 53836 8000
rect 53876 7960 54220 8000
rect 54260 7960 54269 8000
rect 58147 7960 58156 8000
rect 58196 7960 58828 8000
rect 58868 7960 59020 8000
rect 59060 7960 59069 8000
rect 63811 7960 63820 8000
rect 63860 7960 63869 8000
rect 64387 7960 64396 8000
rect 64436 7960 64780 8000
rect 64820 7960 65068 8000
rect 65108 7960 65117 8000
rect 65539 7960 65548 8000
rect 65588 7960 66316 8000
rect 66356 7960 66365 8000
rect 73507 7960 73516 8000
rect 73556 7960 75532 8000
rect 75572 7960 75581 8000
rect 76099 7960 76108 8000
rect 76148 7960 76157 8000
rect 77251 7960 77260 8000
rect 77300 7960 78028 8000
rect 78068 7960 78077 8000
rect 53260 7832 53300 7960
rect 63820 7916 63860 7960
rect 66307 7959 66365 7960
rect 76108 7916 76148 7960
rect 63820 7876 65260 7916
rect 65300 7876 65740 7916
rect 65780 7876 65789 7916
rect 75619 7876 75628 7916
rect 75668 7876 76148 7916
rect 2563 7792 2572 7832
rect 2612 7792 2764 7832
rect 2804 7792 2813 7832
rect 44419 7792 44428 7832
rect 44468 7792 44812 7832
rect 44852 7792 44861 7832
rect 44908 7792 46828 7832
rect 46868 7792 47884 7832
rect 47924 7792 47933 7832
rect 48739 7792 48748 7832
rect 48788 7792 48797 7832
rect 52963 7792 52972 7832
rect 53012 7792 53300 7832
rect 60355 7792 60364 7832
rect 60404 7792 64684 7832
rect 64724 7792 65644 7832
rect 65684 7792 65693 7832
rect 75715 7792 75724 7832
rect 75764 7792 76012 7832
rect 76052 7792 76061 7832
rect 44908 7748 44948 7792
rect 47884 7748 47924 7792
rect 3715 7708 3724 7748
rect 3764 7708 5164 7748
rect 5204 7708 7468 7748
rect 7508 7708 7517 7748
rect 43267 7708 43276 7748
rect 43316 7708 44236 7748
rect 44276 7708 44948 7748
rect 45379 7708 45388 7748
rect 45428 7708 47500 7748
rect 47540 7708 47549 7748
rect 47884 7708 49708 7748
rect 49748 7708 49757 7748
rect 60163 7708 60172 7748
rect 60212 7708 60556 7748
rect 60596 7708 60605 7748
rect 62179 7708 62188 7748
rect 62228 7708 63628 7748
rect 63668 7708 63677 7748
rect 65155 7708 65164 7748
rect 65204 7708 66028 7748
rect 66068 7708 68428 7748
rect 68468 7708 68477 7748
rect 70339 7708 70348 7748
rect 70388 7708 71020 7748
rect 71060 7708 71069 7748
rect 48835 7664 48893 7665
rect 48835 7624 48844 7664
rect 48884 7624 49036 7664
rect 49076 7624 49085 7664
rect 48835 7623 48893 7624
rect 1027 7540 1036 7580
rect 1076 7540 1804 7580
rect 1844 7540 1853 7580
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 15103 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 15489 7580
rect 27103 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 27489 7580
rect 39103 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 39489 7580
rect 51103 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 51489 7580
rect 63103 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 63489 7580
rect 75103 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 75489 7580
rect 76195 7412 76253 7413
rect 47491 7372 47500 7412
rect 47540 7372 47788 7412
rect 47828 7372 47980 7412
rect 48020 7372 48364 7412
rect 48404 7372 48413 7412
rect 76110 7372 76204 7412
rect 76244 7372 76253 7412
rect 76195 7371 76253 7372
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 75811 7288 75820 7328
rect 75860 7288 75900 7328
rect 77347 7288 77356 7328
rect 77396 7288 77836 7328
rect 77876 7288 77885 7328
rect 0 7268 80 7288
rect 75820 7244 75860 7288
rect 50467 7204 50476 7244
rect 50516 7204 52876 7244
rect 52916 7204 52925 7244
rect 53443 7204 53452 7244
rect 53492 7204 53740 7244
rect 53780 7204 54700 7244
rect 54740 7204 54749 7244
rect 59683 7204 59692 7244
rect 59732 7204 60460 7244
rect 60500 7204 60509 7244
rect 69859 7204 69868 7244
rect 69908 7204 70348 7244
rect 70388 7204 70397 7244
rect 75427 7204 75436 7244
rect 75476 7204 76204 7244
rect 76244 7204 76253 7244
rect 76579 7204 76588 7244
rect 76628 7204 77164 7244
rect 77204 7204 77213 7244
rect 77635 7160 77693 7161
rect 2947 7120 2956 7160
rect 2996 7120 4972 7160
rect 5012 7120 5021 7160
rect 53059 7120 53068 7160
rect 53108 7120 53300 7160
rect 58915 7120 58924 7160
rect 58964 7120 60844 7160
rect 60884 7120 61036 7160
rect 61076 7120 61085 7160
rect 64099 7120 64108 7160
rect 64148 7120 64300 7160
rect 64340 7120 64349 7160
rect 64963 7120 64972 7160
rect 65012 7120 65740 7160
rect 65780 7120 65836 7160
rect 65876 7120 66604 7160
rect 66644 7120 66653 7160
rect 67843 7120 67852 7160
rect 67892 7120 68140 7160
rect 68180 7120 69964 7160
rect 70004 7120 70013 7160
rect 70147 7120 70156 7160
rect 70196 7120 70540 7160
rect 70580 7120 70589 7160
rect 71971 7120 71980 7160
rect 72020 7120 72652 7160
rect 72692 7120 72701 7160
rect 75715 7120 75724 7160
rect 75764 7120 76684 7160
rect 76724 7120 77260 7160
rect 77300 7120 77309 7160
rect 77550 7120 77644 7160
rect 77684 7120 77693 7160
rect 53260 7076 53300 7120
rect 77635 7119 77693 7120
rect 2275 7036 2284 7076
rect 2324 7036 4300 7076
rect 4340 7036 4780 7076
rect 4820 7036 4829 7076
rect 53260 7036 53356 7076
rect 53396 7036 53405 7076
rect 59203 7036 59212 7076
rect 59252 7036 60076 7076
rect 60116 7036 60125 7076
rect 63907 7036 63916 7076
rect 63956 7036 64876 7076
rect 64916 7036 64925 7076
rect 66787 7036 66796 7076
rect 66836 7036 69100 7076
rect 69140 7036 69149 7076
rect 75811 7036 75820 7076
rect 75860 7036 76108 7076
rect 76148 7036 76157 7076
rect 65251 6868 65260 6908
rect 65300 6868 65548 6908
rect 65588 6868 66220 6908
rect 66260 6868 66269 6908
rect 76195 6824 76253 6825
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 16343 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 16729 6824
rect 28343 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 28729 6824
rect 40343 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 40729 6824
rect 52343 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 52729 6824
rect 57763 6784 57772 6824
rect 57812 6784 59020 6824
rect 59060 6784 59732 6824
rect 64343 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 64729 6824
rect 71779 6784 71788 6824
rect 71828 6784 71980 6824
rect 72020 6784 72029 6824
rect 75811 6784 75820 6824
rect 75860 6784 76204 6824
rect 76244 6784 76253 6824
rect 76343 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 76729 6824
rect 59692 6740 59732 6784
rect 76195 6783 76253 6784
rect 59683 6700 59692 6740
rect 59732 6700 63916 6740
rect 63956 6700 64780 6740
rect 64820 6700 64829 6740
rect 1507 6616 1516 6656
rect 1556 6616 2188 6656
rect 2228 6616 2237 6656
rect 58339 6616 58348 6656
rect 58388 6616 58828 6656
rect 58868 6616 58877 6656
rect 59011 6616 59020 6656
rect 59060 6616 63380 6656
rect 3619 6532 3628 6572
rect 3668 6532 3916 6572
rect 3956 6532 4204 6572
rect 4244 6532 7468 6572
rect 7508 6532 7517 6572
rect 54211 6532 54220 6572
rect 54260 6532 54604 6572
rect 54644 6532 54653 6572
rect 59500 6532 59692 6572
rect 59732 6532 59741 6572
rect 0 6488 80 6508
rect 59500 6488 59540 6532
rect 63340 6488 63380 6616
rect 74851 6532 74860 6572
rect 74900 6532 75724 6572
rect 75764 6532 75773 6572
rect 76483 6532 76492 6572
rect 76532 6532 77644 6572
rect 77684 6532 79468 6572
rect 79508 6532 79517 6572
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 3523 6448 3532 6488
rect 3572 6448 4492 6488
rect 4532 6448 4541 6488
rect 50083 6448 50092 6488
rect 50132 6448 50860 6488
rect 50900 6448 51724 6488
rect 51764 6448 51773 6488
rect 54403 6448 54412 6488
rect 54452 6448 54796 6488
rect 54836 6448 54845 6488
rect 58051 6448 58060 6488
rect 58100 6448 58540 6488
rect 58580 6448 58589 6488
rect 58819 6448 58828 6488
rect 58868 6448 59212 6488
rect 59252 6448 59261 6488
rect 59491 6448 59500 6488
rect 59540 6448 59549 6488
rect 59779 6448 59788 6488
rect 59828 6448 60172 6488
rect 60212 6448 60221 6488
rect 61315 6448 61324 6488
rect 61364 6448 61900 6488
rect 61940 6448 61949 6488
rect 63340 6448 64108 6488
rect 64148 6448 65260 6488
rect 65300 6448 65309 6488
rect 65923 6448 65932 6488
rect 65972 6448 66796 6488
rect 66836 6448 66845 6488
rect 69955 6448 69964 6488
rect 70004 6448 70444 6488
rect 70484 6448 71884 6488
rect 71924 6448 72940 6488
rect 72980 6448 73228 6488
rect 73268 6448 73277 6488
rect 73603 6448 73612 6488
rect 73652 6448 75628 6488
rect 75668 6448 76300 6488
rect 76340 6448 76588 6488
rect 76628 6448 76637 6488
rect 0 6428 80 6448
rect 45475 6364 45484 6404
rect 45524 6364 47116 6404
rect 47156 6364 47308 6404
rect 47348 6364 47357 6404
rect 57859 6364 57868 6404
rect 57908 6364 58732 6404
rect 58772 6364 59020 6404
rect 59060 6364 59069 6404
rect 2371 6280 2380 6320
rect 2420 6280 2572 6320
rect 2612 6280 2621 6320
rect 45571 6280 45580 6320
rect 45620 6280 47404 6320
rect 47444 6280 47453 6320
rect 56803 6280 56812 6320
rect 56852 6280 58060 6320
rect 58100 6280 58109 6320
rect 58243 6280 58252 6320
rect 58292 6280 60268 6320
rect 60308 6280 60652 6320
rect 60692 6280 60701 6320
rect 65347 6280 65356 6320
rect 65396 6280 65836 6320
rect 65876 6280 65885 6320
rect 74755 6280 74764 6320
rect 74804 6280 75628 6320
rect 75668 6280 75677 6320
rect 48163 6236 48221 6237
rect 7459 6196 7468 6236
rect 7508 6196 48172 6236
rect 48212 6196 48221 6236
rect 51235 6196 51244 6236
rect 51284 6196 51293 6236
rect 51427 6196 51436 6236
rect 51476 6196 52396 6236
rect 52436 6196 52445 6236
rect 63427 6196 63436 6236
rect 63476 6196 63572 6236
rect 48163 6195 48221 6196
rect 51244 6152 51284 6196
rect 50371 6112 50380 6152
rect 50420 6112 60940 6152
rect 60980 6112 60989 6152
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 4195 6028 4204 6068
rect 4244 6028 4972 6068
rect 5012 6028 5021 6068
rect 15103 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 15489 6068
rect 27103 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 27489 6068
rect 39103 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 39489 6068
rect 51103 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 51489 6068
rect 63103 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 63489 6068
rect 63532 5900 63572 6196
rect 69379 6028 69388 6068
rect 69428 6028 69772 6068
rect 69812 6028 69821 6068
rect 75103 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 75489 6068
rect 5059 5860 5068 5900
rect 5108 5860 6316 5900
rect 6356 5860 6365 5900
rect 48547 5860 48556 5900
rect 48596 5860 48748 5900
rect 48788 5860 48797 5900
rect 63331 5860 63340 5900
rect 63380 5860 63572 5900
rect 69187 5860 69196 5900
rect 69236 5860 69772 5900
rect 69812 5860 69821 5900
rect 47395 5776 47404 5816
rect 47444 5776 47596 5816
rect 47636 5776 47645 5816
rect 52771 5776 52780 5816
rect 52820 5776 53164 5816
rect 53204 5776 53213 5816
rect 64195 5776 64204 5816
rect 64244 5776 64253 5816
rect 64579 5776 64588 5816
rect 64628 5776 65068 5816
rect 65108 5776 65117 5816
rect 71971 5776 71980 5816
rect 72020 5776 72212 5816
rect 64204 5732 64244 5776
rect 72172 5732 72212 5776
rect 1507 5692 1516 5732
rect 1556 5692 2956 5732
rect 2996 5692 3628 5732
rect 3668 5692 4108 5732
rect 4148 5692 4157 5732
rect 48451 5692 48460 5732
rect 48500 5692 48509 5732
rect 52675 5692 52684 5732
rect 52724 5692 53548 5732
rect 53588 5692 55852 5732
rect 55892 5692 57388 5732
rect 57428 5692 57964 5732
rect 58004 5692 60076 5732
rect 60116 5692 60125 5732
rect 60643 5692 60652 5732
rect 60692 5692 61996 5732
rect 62036 5692 63628 5732
rect 63668 5692 63677 5732
rect 64204 5692 65164 5732
rect 65204 5692 65213 5732
rect 69292 5692 71692 5732
rect 71732 5692 71741 5732
rect 72163 5692 72172 5732
rect 72212 5692 72221 5732
rect 0 5648 80 5668
rect 48460 5648 48500 5692
rect 69292 5648 69332 5692
rect 71299 5648 71357 5649
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 5731 5608 5740 5648
rect 5780 5608 6220 5648
rect 6260 5608 6269 5648
rect 47395 5608 47404 5648
rect 47444 5608 49132 5648
rect 49172 5608 49181 5648
rect 52291 5608 52300 5648
rect 52340 5608 52349 5648
rect 52963 5608 52972 5648
rect 53012 5608 53932 5648
rect 53972 5608 54220 5648
rect 54260 5608 54269 5648
rect 54691 5608 54700 5648
rect 54740 5608 57004 5648
rect 57044 5608 57053 5648
rect 59395 5608 59404 5648
rect 59444 5608 61324 5648
rect 61364 5608 61373 5648
rect 61507 5608 61516 5648
rect 61556 5608 62476 5648
rect 62516 5608 63532 5648
rect 63572 5608 64204 5648
rect 64244 5608 64253 5648
rect 64771 5608 64780 5648
rect 64820 5608 66220 5648
rect 66260 5608 66508 5648
rect 66548 5608 66557 5648
rect 69091 5608 69100 5648
rect 69140 5608 69292 5648
rect 69332 5608 69341 5648
rect 69955 5608 69964 5648
rect 70004 5608 70013 5648
rect 70819 5608 70828 5648
rect 70868 5608 71308 5648
rect 71348 5608 71357 5648
rect 71587 5608 71596 5648
rect 71636 5608 72748 5648
rect 72788 5608 74380 5648
rect 74420 5608 74429 5648
rect 76387 5608 76396 5648
rect 76436 5608 77260 5648
rect 77300 5608 77309 5648
rect 0 5588 80 5608
rect 52300 5564 52340 5608
rect 1219 5524 1228 5564
rect 1268 5524 2188 5564
rect 2228 5524 2237 5564
rect 48355 5524 48364 5564
rect 48404 5524 50380 5564
rect 50420 5524 50429 5564
rect 52300 5524 54316 5564
rect 54356 5524 54365 5564
rect 54700 5480 54740 5608
rect 69964 5564 70004 5608
rect 71299 5607 71357 5608
rect 54883 5524 54892 5564
rect 54932 5524 56236 5564
rect 56276 5524 58156 5564
rect 58196 5524 58205 5564
rect 63619 5524 63628 5564
rect 63668 5524 67948 5564
rect 67988 5524 67997 5564
rect 69964 5524 71788 5564
rect 71828 5524 72268 5564
rect 72308 5524 72317 5564
rect 66307 5480 66365 5481
rect 1411 5440 1420 5480
rect 1460 5440 1708 5480
rect 1748 5440 1757 5480
rect 47875 5440 47884 5480
rect 47924 5440 48940 5480
rect 48980 5440 48989 5480
rect 54115 5440 54124 5480
rect 54164 5440 54740 5480
rect 58819 5440 58828 5480
rect 58868 5440 59308 5480
rect 59348 5440 59357 5480
rect 62947 5440 62956 5480
rect 62996 5440 64684 5480
rect 64724 5440 64733 5480
rect 65539 5440 65548 5480
rect 65588 5440 66124 5480
rect 66164 5440 66173 5480
rect 66307 5440 66316 5480
rect 66356 5440 66450 5480
rect 76483 5440 76492 5480
rect 76532 5440 76541 5480
rect 66307 5439 66365 5440
rect 76492 5396 76532 5440
rect 64771 5356 64780 5396
rect 64820 5356 65260 5396
rect 65300 5356 65309 5396
rect 76108 5356 76532 5396
rect 76108 5312 76148 5356
rect 3427 5272 3436 5312
rect 3476 5272 4012 5312
rect 4052 5272 4061 5312
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 16343 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 16729 5312
rect 28343 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 28729 5312
rect 40343 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 40729 5312
rect 52343 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 52729 5312
rect 64343 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 64729 5312
rect 76099 5272 76108 5312
rect 76148 5272 76157 5312
rect 76343 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 76729 5312
rect 2860 5188 3532 5228
rect 3572 5188 6124 5228
rect 6164 5188 6173 5228
rect 2860 5144 2900 5188
rect 2275 5104 2284 5144
rect 2324 5104 2900 5144
rect 3907 5104 3916 5144
rect 3956 5104 5932 5144
rect 5972 5104 5981 5144
rect 49123 5104 49132 5144
rect 49172 5104 52012 5144
rect 52052 5104 52300 5144
rect 52340 5104 53300 5144
rect 61027 5104 61036 5144
rect 61076 5104 61420 5144
rect 61460 5104 61469 5144
rect 64867 5104 64876 5144
rect 64916 5104 65644 5144
rect 65684 5104 65693 5144
rect 53260 5060 53300 5104
rect 2755 5020 2764 5060
rect 2804 5020 4300 5060
rect 4340 5020 5740 5060
rect 5780 5020 6508 5060
rect 6548 5020 6557 5060
rect 45667 5020 45676 5060
rect 45716 5020 47308 5060
rect 47348 5020 47357 5060
rect 48547 5020 48556 5060
rect 48596 5020 49228 5060
rect 49268 5020 49277 5060
rect 51811 5020 51820 5060
rect 51860 5020 52588 5060
rect 52628 5020 52637 5060
rect 53251 5020 53260 5060
rect 53300 5020 53309 5060
rect 60163 5020 60172 5060
rect 60212 5020 60460 5060
rect 60500 5020 61612 5060
rect 61652 5020 61661 5060
rect 63340 5020 65164 5060
rect 65204 5020 66124 5060
rect 66164 5020 66173 5060
rect 3427 4936 3436 4976
rect 3476 4936 4684 4976
rect 4724 4936 4733 4976
rect 48259 4936 48268 4976
rect 48308 4936 48460 4976
rect 48500 4936 48509 4976
rect 52099 4936 52108 4976
rect 52148 4936 52492 4976
rect 52532 4936 53452 4976
rect 53492 4936 53501 4976
rect 55939 4936 55948 4976
rect 55988 4936 56332 4976
rect 56372 4936 56381 4976
rect 59203 4936 59212 4976
rect 59252 4936 59692 4976
rect 59732 4936 59741 4976
rect 60067 4936 60076 4976
rect 60116 4936 60940 4976
rect 60980 4936 61516 4976
rect 61556 4936 61565 4976
rect 63340 4892 63380 5020
rect 63619 4936 63628 4976
rect 63668 4936 63916 4976
rect 63956 4936 65548 4976
rect 65588 4936 65597 4976
rect 65731 4936 65740 4976
rect 65780 4936 66508 4976
rect 66548 4936 66557 4976
rect 70819 4936 70828 4976
rect 70868 4936 71500 4976
rect 71540 4936 71549 4976
rect 71875 4936 71884 4976
rect 71924 4936 72172 4976
rect 72212 4936 72221 4976
rect 76579 4936 76588 4976
rect 76628 4936 77356 4976
rect 77396 4936 77405 4976
rect 61603 4852 61612 4892
rect 61652 4852 63380 4892
rect 71308 4852 71788 4892
rect 71828 4852 71837 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 51619 4768 51628 4808
rect 51668 4768 54028 4808
rect 54068 4768 55660 4808
rect 55700 4768 56332 4808
rect 56372 4768 56381 4808
rect 63340 4768 68236 4808
rect 68276 4768 68285 4808
rect 0 4748 80 4768
rect 63340 4724 63380 4768
rect 71308 4724 71348 4852
rect 74467 4768 74476 4808
rect 74516 4768 74860 4808
rect 74900 4768 74909 4808
rect 77443 4768 77452 4808
rect 77492 4768 77836 4808
rect 77876 4768 77885 4808
rect 56419 4684 56428 4724
rect 56468 4684 58540 4724
rect 58580 4684 63380 4724
rect 67747 4684 67756 4724
rect 67796 4684 68812 4724
rect 68852 4684 68861 4724
rect 69187 4684 69196 4724
rect 69236 4684 71308 4724
rect 71348 4684 71357 4724
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 15103 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 15489 4556
rect 27103 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 27489 4556
rect 39103 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 39489 4556
rect 51103 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 51489 4556
rect 63103 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 63489 4556
rect 75103 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 75489 4556
rect 70147 4472 70205 4473
rect 66691 4432 66700 4472
rect 66740 4432 68812 4472
rect 68852 4432 70156 4472
rect 70196 4432 70205 4472
rect 51523 4348 51532 4388
rect 51572 4348 52300 4388
rect 52340 4348 52349 4388
rect 53539 4348 53548 4388
rect 53588 4348 54892 4388
rect 54932 4348 54941 4388
rect 55843 4348 55852 4388
rect 55892 4348 56716 4388
rect 56756 4348 57196 4388
rect 57236 4348 57245 4388
rect 66700 4304 66740 4432
rect 70147 4431 70205 4432
rect 76195 4388 76253 4389
rect 70435 4348 70444 4388
rect 70484 4348 70636 4388
rect 70676 4348 71404 4388
rect 71444 4348 72460 4388
rect 72500 4348 72844 4388
rect 72884 4348 72893 4388
rect 76110 4348 76204 4388
rect 76244 4348 76253 4388
rect 76195 4347 76253 4348
rect 3811 4264 3820 4304
rect 3860 4264 4396 4304
rect 4436 4264 7660 4304
rect 7700 4264 7709 4304
rect 51907 4264 51916 4304
rect 51956 4264 52684 4304
rect 52724 4264 54700 4304
rect 54740 4264 55180 4304
rect 55220 4264 55229 4304
rect 57283 4264 57292 4304
rect 57332 4264 57964 4304
rect 58004 4264 58013 4304
rect 59395 4264 59404 4304
rect 59444 4264 59596 4304
rect 59636 4264 61804 4304
rect 61844 4264 61853 4304
rect 62755 4264 62764 4304
rect 62804 4264 64012 4304
rect 64052 4264 64061 4304
rect 65827 4264 65836 4304
rect 65876 4264 66740 4304
rect 68707 4264 68716 4304
rect 68756 4264 69004 4304
rect 69044 4264 70252 4304
rect 70292 4264 70732 4304
rect 70772 4264 70781 4304
rect 71299 4264 71308 4304
rect 71348 4264 72076 4304
rect 72116 4264 72125 4304
rect 73699 4264 73708 4304
rect 73748 4264 74284 4304
rect 74324 4264 74333 4304
rect 75811 4264 75820 4304
rect 75860 4264 76876 4304
rect 76916 4264 76925 4304
rect 77827 4264 77836 4304
rect 77876 4264 78412 4304
rect 78452 4264 79468 4304
rect 79508 4264 79517 4304
rect 4483 4180 4492 4220
rect 4532 4180 4780 4220
rect 4820 4180 4829 4220
rect 50659 4180 50668 4220
rect 50708 4180 53068 4220
rect 53108 4180 55660 4220
rect 55700 4180 55709 4220
rect 58627 4180 58636 4220
rect 58676 4180 59116 4220
rect 59156 4180 59980 4220
rect 60020 4180 60029 4220
rect 74467 4180 74476 4220
rect 74516 4180 76396 4220
rect 76436 4180 76445 4220
rect 3043 4096 3052 4136
rect 3092 4096 4876 4136
rect 4916 4096 4925 4136
rect 5059 4096 5068 4136
rect 5108 4096 6316 4136
rect 6356 4096 6365 4136
rect 55555 4096 55564 4136
rect 55604 4096 57004 4136
rect 57044 4096 57053 4136
rect 58243 4096 58252 4136
rect 58292 4096 58924 4136
rect 58964 4096 60748 4136
rect 60788 4096 61228 4136
rect 61268 4096 61277 4136
rect 68803 4096 68812 4136
rect 68852 4096 70444 4136
rect 70484 4096 70493 4136
rect 74563 4096 74572 4136
rect 74612 4096 74764 4136
rect 74804 4096 75724 4136
rect 75764 4096 76780 4136
rect 76820 4096 76829 4136
rect 2659 4012 2668 4052
rect 2708 4012 3724 4052
rect 3764 4012 3916 4052
rect 3956 4012 3965 4052
rect 50851 4012 50860 4052
rect 50900 4012 54604 4052
rect 54644 4012 54653 4052
rect 65251 4012 65260 4052
rect 65300 4012 65932 4052
rect 65972 4012 65981 4052
rect 0 3968 80 3988
rect 0 3928 1036 3968
rect 1076 3928 1085 3968
rect 2563 3928 2572 3968
rect 2612 3928 3532 3968
rect 3572 3928 4012 3968
rect 4052 3928 4588 3968
rect 4628 3928 4637 3968
rect 50755 3928 50764 3968
rect 50804 3928 52972 3968
rect 53012 3928 55756 3968
rect 55796 3928 55805 3968
rect 55939 3928 55948 3968
rect 55988 3928 56524 3968
rect 56564 3928 56573 3968
rect 0 3908 80 3928
rect 53827 3844 53836 3884
rect 53876 3844 56140 3884
rect 56180 3844 56189 3884
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 16343 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 16729 3800
rect 28343 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 28729 3800
rect 40343 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 40729 3800
rect 52343 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 52729 3800
rect 55075 3760 55084 3800
rect 55124 3760 55756 3800
rect 55796 3760 55805 3800
rect 64343 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 64729 3800
rect 76343 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 76729 3800
rect 71299 3716 71357 3717
rect 59491 3676 59500 3716
rect 59540 3676 62092 3716
rect 62132 3676 67372 3716
rect 67412 3676 67421 3716
rect 71299 3676 71308 3716
rect 71348 3676 71788 3716
rect 71828 3676 71837 3716
rect 71299 3675 71357 3676
rect 49603 3592 49612 3632
rect 49652 3592 50188 3632
rect 50228 3592 50237 3632
rect 50851 3592 50860 3632
rect 50900 3592 52012 3632
rect 52052 3592 52061 3632
rect 62851 3592 62860 3632
rect 62900 3592 64012 3632
rect 64052 3592 64061 3632
rect 68995 3592 69004 3632
rect 69044 3592 69292 3632
rect 69332 3592 69341 3632
rect 70723 3592 70732 3632
rect 70772 3592 72076 3632
rect 72116 3592 72125 3632
rect 76003 3592 76012 3632
rect 76052 3592 76300 3632
rect 76340 3592 76349 3632
rect 1315 3508 1324 3548
rect 1364 3508 2956 3548
rect 2996 3508 3005 3548
rect 4387 3508 4396 3548
rect 4436 3508 4876 3548
rect 4916 3508 4925 3548
rect 51628 3508 53836 3548
rect 53876 3508 53885 3548
rect 56131 3508 56140 3548
rect 56180 3508 57100 3548
rect 57140 3508 57149 3548
rect 69955 3508 69964 3548
rect 70004 3508 70636 3548
rect 70676 3508 71404 3548
rect 71444 3508 71453 3548
rect 71587 3508 71596 3548
rect 71636 3508 72268 3548
rect 72308 3508 73708 3548
rect 73748 3508 73757 3548
rect 75811 3508 75820 3548
rect 75860 3508 76780 3548
rect 76820 3508 76829 3548
rect 51628 3464 51668 3508
rect 76195 3464 76253 3465
rect 51619 3424 51628 3464
rect 51668 3424 51677 3464
rect 52675 3424 52684 3464
rect 52724 3424 54508 3464
rect 54548 3424 56620 3464
rect 56660 3424 56669 3464
rect 58819 3424 58828 3464
rect 58868 3424 59692 3464
rect 59732 3424 59741 3464
rect 63907 3424 63916 3464
rect 63956 3424 63965 3464
rect 64579 3424 64588 3464
rect 64628 3424 65260 3464
rect 65300 3424 65309 3464
rect 68899 3424 68908 3464
rect 68948 3424 68957 3464
rect 70243 3424 70252 3464
rect 70292 3424 72460 3464
rect 72500 3424 72748 3464
rect 72788 3424 73132 3464
rect 73172 3424 74572 3464
rect 74612 3424 74621 3464
rect 76099 3424 76108 3464
rect 76148 3424 76204 3464
rect 76244 3424 76253 3464
rect 76675 3424 76684 3464
rect 76724 3424 77836 3464
rect 77876 3424 77885 3464
rect 63916 3380 63956 3424
rect 68908 3380 68948 3424
rect 76195 3423 76253 3424
rect 1123 3340 1132 3380
rect 1172 3340 2476 3380
rect 2516 3340 2525 3380
rect 63916 3340 66028 3380
rect 66068 3340 66316 3380
rect 66356 3340 66365 3380
rect 68908 3340 70540 3380
rect 70580 3340 70924 3380
rect 70964 3340 74860 3380
rect 74900 3340 74909 3380
rect 1891 3256 1900 3296
rect 1940 3256 2668 3296
rect 2708 3256 2717 3296
rect 50083 3256 50092 3296
rect 50132 3256 51724 3296
rect 51764 3256 52588 3296
rect 52628 3256 52637 3296
rect 64099 3256 64108 3296
rect 64148 3256 65452 3296
rect 65492 3256 65501 3296
rect 68227 3256 68236 3296
rect 68276 3256 69772 3296
rect 69812 3256 71692 3296
rect 71732 3256 71741 3296
rect 73987 3256 73996 3296
rect 74036 3256 76396 3296
rect 76436 3256 76780 3296
rect 76820 3256 76829 3296
rect 1603 3172 1612 3212
rect 1652 3172 2572 3212
rect 2612 3172 2621 3212
rect 72835 3172 72844 3212
rect 72884 3172 77452 3212
rect 77492 3172 77836 3212
rect 77876 3172 77885 3212
rect 0 3128 80 3148
rect 0 3088 652 3128
rect 692 3088 701 3128
rect 59011 3088 59020 3128
rect 59060 3088 60556 3128
rect 60596 3088 60605 3128
rect 68707 3088 68716 3128
rect 68756 3088 69004 3128
rect 69044 3088 69053 3128
rect 71683 3088 71692 3128
rect 71732 3088 76012 3128
rect 76052 3088 76061 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 15103 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 15489 3044
rect 27103 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 27489 3044
rect 39103 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 39489 3044
rect 51103 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 51489 3044
rect 59395 3004 59404 3044
rect 59444 3004 60364 3044
rect 60404 3004 60413 3044
rect 63103 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 63489 3044
rect 75103 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 75489 3044
rect 59971 2920 59980 2960
rect 60020 2920 62764 2960
rect 62804 2920 62813 2960
rect 74851 2920 74860 2960
rect 74900 2920 76108 2960
rect 76148 2920 76157 2960
rect 76867 2920 76876 2960
rect 76916 2920 78124 2960
rect 78164 2920 78316 2960
rect 78356 2920 78365 2960
rect 58915 2836 58924 2876
rect 58964 2836 64204 2876
rect 64244 2836 66124 2876
rect 66164 2836 66173 2876
rect 71203 2836 71212 2876
rect 71252 2836 72940 2876
rect 72980 2836 72989 2876
rect 53731 2752 53740 2792
rect 53780 2752 55756 2792
rect 55796 2752 55805 2792
rect 56227 2752 56236 2792
rect 56276 2752 56524 2792
rect 56564 2752 56908 2792
rect 56948 2752 56957 2792
rect 71875 2752 71884 2792
rect 71924 2752 73612 2792
rect 73652 2752 73661 2792
rect 73891 2752 73900 2792
rect 73940 2752 74668 2792
rect 74708 2752 74717 2792
rect 1699 2668 1708 2708
rect 1748 2668 3380 2708
rect 55843 2668 55852 2708
rect 55892 2668 57292 2708
rect 57332 2668 57341 2708
rect 58723 2668 58732 2708
rect 58772 2668 59020 2708
rect 59060 2668 60364 2708
rect 60404 2668 60413 2708
rect 64483 2668 64492 2708
rect 64532 2668 64780 2708
rect 64820 2668 64829 2708
rect 71011 2668 71020 2708
rect 71060 2668 71308 2708
rect 71348 2668 71357 2708
rect 71779 2668 71788 2708
rect 71828 2668 72076 2708
rect 72116 2668 72125 2708
rect 72931 2668 72940 2708
rect 72980 2668 74188 2708
rect 74228 2668 74237 2708
rect 74467 2668 74476 2708
rect 74516 2668 76396 2708
rect 76436 2668 77356 2708
rect 77396 2668 77405 2708
rect 3340 2624 3380 2668
rect 51715 2624 51773 2625
rect 75715 2624 75773 2625
rect 77347 2624 77405 2625
rect 2371 2584 2380 2624
rect 2420 2584 3052 2624
rect 3092 2584 3101 2624
rect 3331 2584 3340 2624
rect 3380 2584 6028 2624
rect 6068 2584 6077 2624
rect 51715 2584 51724 2624
rect 51764 2584 72172 2624
rect 72212 2584 72221 2624
rect 73699 2584 73708 2624
rect 73748 2584 74284 2624
rect 74324 2584 74764 2624
rect 74804 2584 75724 2624
rect 75764 2584 75773 2624
rect 77059 2584 77068 2624
rect 77108 2584 77356 2624
rect 77396 2584 78892 2624
rect 78932 2584 78941 2624
rect 51715 2583 51773 2584
rect 75715 2583 75773 2584
rect 77347 2583 77405 2584
rect 71299 2540 71357 2541
rect 53155 2500 53164 2540
rect 53204 2500 56044 2540
rect 56084 2500 57580 2540
rect 57620 2500 57629 2540
rect 59779 2500 59788 2540
rect 59828 2500 60652 2540
rect 60692 2500 61612 2540
rect 61652 2500 61661 2540
rect 64387 2500 64396 2540
rect 64436 2500 64780 2540
rect 64820 2500 64829 2540
rect 68323 2500 68332 2540
rect 68372 2500 69868 2540
rect 69908 2500 70580 2540
rect 70540 2456 70580 2500
rect 71299 2500 71308 2540
rect 71348 2500 73996 2540
rect 74036 2500 74045 2540
rect 71299 2499 71357 2500
rect 63811 2416 63820 2456
rect 63860 2416 64684 2456
rect 64724 2416 65740 2456
rect 65780 2416 65789 2456
rect 67363 2416 67372 2456
rect 67412 2416 68140 2456
rect 68180 2416 68189 2456
rect 70540 2416 72076 2456
rect 72116 2416 75820 2456
rect 75860 2416 76108 2456
rect 76148 2416 76157 2456
rect 76771 2416 76780 2456
rect 76820 2416 77164 2456
rect 77204 2416 77213 2456
rect 77347 2416 77356 2456
rect 77396 2416 78700 2456
rect 78740 2416 78749 2456
rect 68227 2332 68236 2372
rect 68276 2332 69196 2372
rect 69236 2332 71020 2372
rect 71060 2332 71212 2372
rect 71252 2332 71261 2372
rect 0 2288 80 2308
rect 71299 2288 71357 2289
rect 0 2248 1036 2288
rect 1076 2248 1085 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 16343 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 16729 2288
rect 28343 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 28729 2288
rect 40343 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 40729 2288
rect 52343 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 52729 2288
rect 64343 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 64729 2288
rect 67939 2248 67948 2288
rect 67988 2248 71308 2288
rect 71348 2248 71357 2288
rect 74467 2248 74476 2288
rect 74516 2248 74668 2288
rect 74708 2248 74717 2288
rect 76343 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 76729 2288
rect 0 2228 80 2248
rect 71299 2247 71357 2248
rect 55459 2164 55468 2204
rect 55508 2164 56044 2204
rect 56084 2164 56093 2204
rect 73987 2164 73996 2204
rect 74036 2164 76972 2204
rect 77012 2164 78220 2204
rect 78260 2164 78269 2204
rect 55843 2080 55852 2120
rect 55892 2080 56524 2120
rect 56564 2080 57196 2120
rect 57236 2080 57245 2120
rect 65155 2080 65164 2120
rect 65204 2080 66892 2120
rect 66932 2080 66941 2120
rect 55939 1912 55948 1952
rect 55988 1912 56332 1952
rect 56372 1912 56381 1952
rect 56995 1912 57004 1952
rect 57044 1912 57388 1952
rect 57428 1912 57437 1952
rect 57859 1912 57868 1952
rect 57908 1912 59116 1952
rect 59156 1912 60460 1952
rect 60500 1912 60940 1952
rect 60980 1912 60989 1952
rect 63043 1912 63052 1952
rect 63092 1912 65740 1952
rect 65780 1912 67276 1952
rect 67316 1912 67468 1952
rect 67508 1912 70060 1952
rect 70100 1912 70252 1952
rect 70292 1912 70301 1952
rect 70915 1912 70924 1952
rect 70964 1912 71788 1952
rect 71828 1912 71837 1952
rect 73795 1912 73804 1952
rect 73844 1912 74572 1952
rect 74612 1912 74621 1952
rect 75235 1912 75244 1952
rect 75284 1912 77740 1952
rect 77780 1912 78412 1952
rect 78452 1912 78461 1952
rect 67555 1828 67564 1868
rect 67604 1828 68524 1868
rect 68564 1828 68573 1868
rect 68995 1828 69004 1868
rect 69044 1828 70828 1868
rect 70868 1828 73996 1868
rect 74036 1828 74045 1868
rect 53443 1744 53452 1784
rect 53492 1744 55948 1784
rect 55988 1744 55997 1784
rect 59011 1660 59020 1700
rect 59060 1660 68044 1700
rect 68084 1660 68093 1700
rect 74755 1576 74764 1616
rect 74804 1576 75628 1616
rect 75668 1576 75677 1616
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 15103 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 15489 1532
rect 27103 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 27489 1532
rect 39103 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 39489 1532
rect 51103 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 51489 1532
rect 63103 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 63489 1532
rect 75103 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 75489 1532
rect 57187 1408 57196 1448
rect 57236 1408 59020 1448
rect 59060 1408 59069 1448
rect 64099 1408 64108 1448
rect 64148 1408 65164 1448
rect 65204 1408 65213 1448
rect 58915 1324 58924 1364
rect 58964 1324 59212 1364
rect 59252 1324 59261 1364
rect 61795 1324 61804 1364
rect 61844 1324 62476 1364
rect 62516 1324 62525 1364
rect 59587 1240 59596 1280
rect 59636 1240 60844 1280
rect 60884 1240 60893 1280
rect 62275 1240 62284 1280
rect 62324 1240 64780 1280
rect 64820 1240 64829 1280
rect 78211 1240 78220 1280
rect 78260 1240 79468 1280
rect 79508 1240 79517 1280
rect 55747 1156 55756 1196
rect 55796 1156 56524 1196
rect 56564 1156 56573 1196
rect 60547 1156 60556 1196
rect 60596 1156 62860 1196
rect 62900 1156 62909 1196
rect 66019 1156 66028 1196
rect 66068 1156 67372 1196
rect 67412 1156 67421 1196
rect 56419 1072 56428 1112
rect 56468 1072 57196 1112
rect 57236 1072 57245 1112
rect 57475 1072 57484 1112
rect 57524 1072 58636 1112
rect 58676 1072 58685 1112
rect 59875 1072 59884 1112
rect 59924 1072 60076 1112
rect 60116 1072 70732 1112
rect 70772 1072 71212 1112
rect 71252 1072 71261 1112
rect 73219 1072 73228 1112
rect 73268 1072 73996 1112
rect 74036 1072 74045 1112
rect 76195 1072 76204 1112
rect 76244 1072 76780 1112
rect 76820 1072 78028 1112
rect 78068 1072 78077 1112
rect 61987 988 61996 1028
rect 62036 988 63628 1028
rect 63668 988 63677 1028
rect 58915 904 58924 944
rect 58964 904 60364 944
rect 60404 904 60413 944
rect 62947 904 62956 944
rect 62996 904 63724 944
rect 63764 904 64204 944
rect 64244 904 64253 944
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 16343 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 16729 776
rect 28343 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 28729 776
rect 40343 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 40729 776
rect 52343 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 52729 776
rect 64343 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 64729 776
rect 76343 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 76729 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 59404 38200 59444 38240
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 72460 37360 72500 37400
rect 76972 37360 77012 37400
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 69100 36856 69140 36896
rect 69100 36436 69140 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67564 36268 67604 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 76876 36184 76916 36224
rect 50860 35848 50900 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 67564 33916 67604 33956
rect 76876 33748 76916 33788
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 50860 32824 50900 32864
rect 70636 32572 70676 32612
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 76876 32236 76916 32276
rect 77452 32152 77492 32192
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 51628 31396 51668 31436
rect 71980 31396 72020 31436
rect 77260 31228 77300 31268
rect 71116 31144 71156 31184
rect 76876 31144 76916 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 41164 30556 41204 30596
rect 71980 30556 72020 30596
rect 77260 30556 77300 30596
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 72460 30220 72500 30260
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 76108 30220 76148 30260
rect 77260 30220 77300 30260
rect 40780 30052 40820 30092
rect 71308 30136 71348 30176
rect 71116 29968 71156 30008
rect 71308 29716 71348 29756
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 64012 29128 64052 29168
rect 71404 28792 71444 28832
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 77836 28708 77876 28748
rect 50476 28540 50516 28580
rect 54604 28540 54644 28580
rect 59404 28540 59444 28580
rect 64012 28456 64052 28496
rect 65164 28456 65204 28496
rect 46636 28288 46676 28328
rect 60172 28288 60212 28328
rect 50668 28120 50708 28160
rect 52108 28036 52148 28076
rect 71692 28036 71732 28076
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 52780 27952 52820 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 58252 27616 58292 27656
rect 41068 27532 41108 27572
rect 46348 27532 46388 27572
rect 52012 27448 52052 27488
rect 52780 27448 52820 27488
rect 43084 27364 43124 27404
rect 50764 27364 50804 27404
rect 67564 27532 67604 27572
rect 60172 27364 60212 27404
rect 71980 27448 72020 27488
rect 65164 27280 65204 27320
rect 71404 27280 71444 27320
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 40204 27112 40244 27152
rect 52972 27112 53012 27152
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 58540 27028 58580 27068
rect 50476 26944 50516 26984
rect 50668 26944 50708 26984
rect 40780 26860 40820 26900
rect 58348 26860 58388 26900
rect 60364 26860 60404 26900
rect 40012 26776 40052 26816
rect 41164 26692 41204 26732
rect 53068 26524 53108 26564
rect 71980 26524 72020 26564
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 54508 26440 54548 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 38956 26272 38996 26312
rect 64012 26272 64052 26312
rect 52204 26104 52244 26144
rect 59404 26104 59444 26144
rect 38860 26020 38900 26060
rect 40876 26020 40916 26060
rect 46828 25936 46868 25976
rect 59404 25852 59444 25892
rect 60364 26020 60404 26060
rect 60556 26020 60596 26060
rect 77836 25852 77876 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 41164 25684 41204 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 63916 25600 63956 25640
rect 41068 25516 41108 25556
rect 46156 25264 46196 25304
rect 46636 25264 46676 25304
rect 50668 25264 50708 25304
rect 51628 25180 51668 25220
rect 40012 25096 40052 25136
rect 60364 25096 60404 25136
rect 63916 25012 63956 25052
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 46828 24592 46868 24632
rect 47308 24760 47348 24800
rect 63916 24676 63956 24716
rect 38956 24508 38996 24548
rect 39724 24424 39764 24464
rect 47308 24256 47348 24296
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 51340 23920 51380 23960
rect 54796 23752 54836 23792
rect 55852 23752 55892 23792
rect 56812 23752 56852 23792
rect 57292 23752 57332 23792
rect 70636 23752 70676 23792
rect 71692 23752 71732 23792
rect 76108 23752 76148 23792
rect 76972 23752 77012 23792
rect 77452 23752 77492 23792
rect 79084 23752 79124 23792
rect 51724 23668 51764 23708
rect 46156 23584 46196 23624
rect 58252 23584 58292 23624
rect 60556 23584 60596 23624
rect 56140 23500 56180 23540
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 54796 23416 54836 23456
rect 56812 23416 56852 23456
rect 52492 23248 52532 23288
rect 56812 23248 56852 23288
rect 55660 23164 55700 23204
rect 46060 23080 46100 23120
rect 51340 23080 51380 23120
rect 56140 22996 56180 23036
rect 54700 22828 54740 22868
rect 54412 22744 54452 22784
rect 57676 22744 57695 22784
rect 57695 22744 57716 22784
rect 60556 22744 60596 22784
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 46156 22660 46196 22700
rect 51820 22576 51860 22616
rect 38860 22156 38900 22196
rect 52300 22156 52340 22196
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 38860 21820 38900 21860
rect 52588 21568 52628 21608
rect 51628 21232 51668 21272
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 40204 21064 40244 21104
rect 52300 20896 52340 20936
rect 43084 20812 43124 20852
rect 46060 20812 46100 20852
rect 40204 20728 40244 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 52492 20224 52532 20264
rect 47692 19804 47732 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 11692 19468 11732 19508
rect 40876 19468 40916 19508
rect 40204 19300 40244 19340
rect 39724 19216 39764 19256
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 47404 18880 47444 18920
rect 33292 18796 33332 18836
rect 33484 18544 33524 18584
rect 49036 18712 49076 18752
rect 46156 18544 46196 18584
rect 51916 18544 51956 18584
rect 43084 18460 43124 18500
rect 47404 18460 47444 18500
rect 51820 18460 51860 18500
rect 33484 18376 33524 18416
rect 46252 18376 46292 18416
rect 47692 18376 47732 18416
rect 51340 18376 51380 18416
rect 33292 18292 33332 18332
rect 35404 18292 35444 18332
rect 40204 18208 40244 18248
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 26476 18124 26516 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 26476 17872 26516 17912
rect 26476 17704 26516 17744
rect 25516 17620 25556 17660
rect 46732 17536 46772 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 32812 17284 32852 17324
rect 54316 17200 54345 17240
rect 54345 17200 54356 17240
rect 55084 17200 55124 17240
rect 58252 17200 58292 17240
rect 40876 17116 40916 17156
rect 52300 17116 52340 17156
rect 57868 17116 57908 17156
rect 52588 17032 52628 17072
rect 52780 17032 52820 17072
rect 75724 17200 75764 17240
rect 54700 17032 54740 17072
rect 46156 16948 46196 16988
rect 36652 16864 36692 16904
rect 27532 16780 27572 16820
rect 29644 16780 29684 16820
rect 39724 16780 39764 16820
rect 49036 16780 49076 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 61708 16276 61748 16316
rect 27532 16192 27572 16232
rect 46252 16192 46292 16232
rect 52780 16192 52820 16232
rect 55084 16192 55124 16232
rect 58540 16192 58580 16232
rect 64972 16192 65012 16232
rect 70156 16192 70196 16232
rect 75724 16192 75764 16232
rect 77644 16192 77684 16232
rect 78892 16192 78932 16232
rect 68524 16024 68564 16064
rect 69100 16024 69140 16064
rect 77356 16024 77396 16064
rect 51916 15940 51956 15980
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 60652 15772 60692 15812
rect 47692 15688 47732 15728
rect 33100 15604 33140 15644
rect 47980 15520 48020 15560
rect 4780 15352 4820 15392
rect 33196 15352 33236 15392
rect 62956 15352 62996 15392
rect 63340 15352 63380 15392
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 60748 15016 60788 15056
rect 46732 14764 46772 14804
rect 47980 14764 48020 14804
rect 61900 14848 61940 14888
rect 50764 14764 50804 14804
rect 67180 14764 67220 14804
rect 60748 14680 60788 14720
rect 32332 14512 32372 14552
rect 4876 14428 4916 14468
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 49324 14596 49364 14636
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 52780 14092 52820 14132
rect 1996 14008 2036 14048
rect 57772 14008 57812 14048
rect 63916 13924 63956 13964
rect 69196 13840 69236 13880
rect 68524 13756 68564 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 36652 13420 36692 13460
rect 47692 13420 47732 13460
rect 74860 13420 74900 13460
rect 47980 13252 48020 13292
rect 49324 13168 49364 13208
rect 76204 13168 76244 13208
rect 74860 13084 74900 13124
rect 36364 13000 36404 13040
rect 57868 13000 57908 13040
rect 68908 13000 68948 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 51916 12832 51956 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 2092 12580 2132 12620
rect 4780 12496 4820 12536
rect 63532 12496 63572 12536
rect 63916 12496 63956 12536
rect 36364 12412 36404 12452
rect 1996 12160 2036 12200
rect 51532 12328 51572 12368
rect 36652 12160 36692 12200
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 52204 11908 52244 11948
rect 60652 11908 60692 11948
rect 2092 11824 2132 11864
rect 47692 11740 47732 11780
rect 68908 11656 68948 11696
rect 70540 11572 70580 11612
rect 76396 11572 76436 11612
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 74860 11320 74900 11360
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 4780 11152 4820 11192
rect 4876 10984 4916 11024
rect 40876 10984 40916 11024
rect 49324 10984 49364 11024
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 63532 10396 63572 10436
rect 58924 10228 58964 10268
rect 4780 9976 4820 10016
rect 69100 10060 69140 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 48652 9724 48692 9764
rect 76204 9556 76244 9596
rect 4780 9304 4820 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 50860 8464 50900 8504
rect 76204 8380 76244 8420
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 48844 8296 48884 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 4780 7960 4820 8000
rect 66316 7960 66356 8000
rect 48844 7624 48884 7664
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 76204 7372 76244 7412
rect 77644 7120 77684 7160
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 76204 6784 76244 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 48172 6196 48212 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 71308 5608 71348 5648
rect 66316 5440 66356 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 70156 4432 70196 4472
rect 76204 4348 76244 4388
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 71308 3676 71348 3716
rect 76204 3424 76244 3464
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 51724 2584 51764 2624
rect 75724 2584 75764 2624
rect 77356 2584 77396 2624
rect 71308 2500 71348 2540
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 71308 2248 71348 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 59404 38240 59444 38249
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 50860 35888 50900 35897
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 50860 32864 50900 35848
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 50860 32815 50900 32824
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 51628 31436 51668 31445
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 41164 30596 41204 30605
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 40780 30092 40820 30101
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 40204 27152 40244 27161
rect 40012 26816 40052 26825
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 38956 26312 38996 26321
rect 38860 26060 38900 26071
rect 38860 25985 38900 26020
rect 38859 25976 38901 25985
rect 38859 25936 38860 25976
rect 38900 25936 38901 25976
rect 38859 25927 38901 25936
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 11691 23204 11733 23213
rect 11691 23164 11692 23204
rect 11732 23164 11733 23204
rect 11691 23155 11733 23164
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 11692 19508 11732 23155
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 38860 22196 38900 25927
rect 38956 24548 38996 26272
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 40012 25136 40052 26776
rect 40012 25087 40052 25096
rect 38956 24499 38996 24508
rect 39724 24464 39764 24473
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 38860 21860 38900 22156
rect 38860 21811 38900 21820
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 11692 19459 11732 19468
rect 39724 19256 39764 24424
rect 40204 21104 40244 27112
rect 40780 26900 40820 30052
rect 40780 26851 40820 26860
rect 41068 27572 41108 27581
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 40875 26060 40917 26069
rect 40875 26020 40876 26060
rect 40916 26020 40917 26060
rect 40875 26011 40917 26020
rect 40876 25926 40916 26011
rect 41068 25556 41108 27532
rect 41164 26732 41204 30556
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 50476 28580 50516 28589
rect 46636 28328 46676 28337
rect 46348 27572 46388 27581
rect 46636 27572 46676 28288
rect 46388 27532 46676 27572
rect 46348 27523 46388 27532
rect 41164 25724 41204 26692
rect 41164 25675 41204 25684
rect 43084 27404 43124 27413
rect 43084 26144 43124 27364
rect 43179 26144 43221 26153
rect 43084 26104 43180 26144
rect 43220 26104 43221 26144
rect 41068 25507 41108 25516
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 40204 20768 40244 21064
rect 43084 20852 43124 26104
rect 43179 26095 43221 26104
rect 43180 26076 43220 26095
rect 46156 25304 46196 25313
rect 46156 23624 46196 25264
rect 46636 25304 46676 27532
rect 50476 26984 50516 28540
rect 50476 26935 50516 26944
rect 50668 28160 50708 28169
rect 50668 26984 50708 28120
rect 46636 25255 46676 25264
rect 46828 25976 46868 25985
rect 46828 24632 46868 25936
rect 50668 25304 50708 26944
rect 50668 25255 50708 25264
rect 50764 27404 50804 27413
rect 46828 24583 46868 24592
rect 47308 24800 47348 24809
rect 47308 24296 47348 24760
rect 47308 24247 47348 24256
rect 48171 23708 48213 23717
rect 48171 23668 48172 23708
rect 48212 23668 48213 23708
rect 48171 23659 48213 23668
rect 43084 20803 43124 20812
rect 46060 23120 46100 23129
rect 46060 20852 46100 23080
rect 46156 22700 46196 23584
rect 46156 22651 46196 22660
rect 46060 20803 46100 20812
rect 40204 20719 40244 20728
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 47692 19844 47732 19853
rect 40876 19508 40916 19517
rect 39724 19207 39764 19216
rect 40204 19340 40244 19349
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 33292 18836 33332 18845
rect 33292 18332 33332 18796
rect 33484 18584 33524 18593
rect 33484 18416 33524 18544
rect 33484 18367 33524 18376
rect 33292 18283 33332 18292
rect 35403 18332 35445 18341
rect 35403 18292 35404 18332
rect 35444 18292 35445 18332
rect 35403 18283 35445 18292
rect 35404 18198 35444 18283
rect 40204 18248 40244 19300
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 40204 18199 40244 18208
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 26476 18164 26516 18173
rect 26476 17912 26516 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 26476 17744 26516 17872
rect 26476 17695 26516 17704
rect 25516 17660 25556 17671
rect 25516 17585 25556 17620
rect 25515 17576 25557 17585
rect 25515 17536 25516 17576
rect 25556 17536 25557 17576
rect 25515 17527 25557 17536
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 32812 17324 32852 17333
rect 32812 16997 32852 17284
rect 40876 17156 40916 19468
rect 47404 18920 47444 18929
rect 46156 18584 46196 18593
rect 43083 18500 43125 18509
rect 43083 18460 43084 18500
rect 43124 18460 43125 18500
rect 43083 18451 43125 18460
rect 43084 18366 43124 18451
rect 32811 16988 32853 16997
rect 32811 16948 32812 16988
rect 32852 16948 32853 16988
rect 32811 16939 32853 16948
rect 36651 16904 36693 16913
rect 36651 16864 36652 16904
rect 36692 16864 36693 16904
rect 36651 16855 36693 16864
rect 27532 16820 27572 16829
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 27532 16232 27572 16780
rect 29643 16820 29685 16829
rect 29643 16780 29644 16820
rect 29684 16780 29685 16820
rect 29643 16771 29685 16780
rect 29644 16686 29684 16771
rect 36652 16770 36692 16855
rect 39724 16820 39764 16831
rect 39724 16745 39764 16780
rect 39723 16736 39765 16745
rect 39723 16696 39724 16736
rect 39764 16696 39765 16736
rect 39723 16687 39765 16696
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 27532 16183 27572 16192
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 33100 15644 33140 15653
rect 33140 15604 33236 15644
rect 33100 15595 33140 15604
rect 4780 15392 4820 15401
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 1996 14048 2036 14057
rect 1996 12200 2036 14008
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 1996 12151 2036 12160
rect 2092 12620 2132 12629
rect 2092 11864 2132 12580
rect 4780 12536 4820 15352
rect 33196 15392 33236 15604
rect 33196 15343 33236 15352
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 32331 14552 32373 14561
rect 32331 14512 32332 14552
rect 32372 14512 32373 14552
rect 32331 14503 32373 14512
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 2092 11815 2132 11824
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4780 11192 4820 12496
rect 4780 11143 4820 11152
rect 4876 14468 4916 14477
rect 4876 11024 4916 14428
rect 32332 14418 32372 14503
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 36652 13460 36692 13469
rect 36364 13040 36404 13049
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 36364 12452 36404 13000
rect 36364 12403 36404 12412
rect 36652 12200 36692 13420
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 36652 12151 36692 12160
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 4876 10975 4916 10984
rect 40876 11024 40916 17116
rect 46156 16988 46196 18544
rect 47404 18500 47444 18880
rect 47404 18451 47444 18460
rect 46156 16939 46196 16948
rect 46252 18416 46292 18425
rect 46252 16232 46292 18376
rect 47692 18416 47732 19804
rect 46252 16183 46292 16192
rect 46732 17576 46772 17585
rect 46732 14804 46772 17536
rect 46732 14755 46772 14764
rect 47692 15728 47732 18376
rect 47692 13460 47732 15688
rect 47692 11780 47732 13420
rect 47980 15560 48020 15569
rect 47980 14804 48020 15520
rect 47980 13292 48020 14764
rect 47980 13243 48020 13252
rect 47692 11731 47732 11740
rect 40876 10975 40916 10984
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 4780 10016 4820 10025
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4780 9344 4820 9976
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4780 8000 4820 9304
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 4780 7951 4820 7960
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 48172 6236 48212 23659
rect 48651 23624 48693 23633
rect 48651 23584 48652 23624
rect 48692 23584 48693 23624
rect 48651 23575 48693 23584
rect 48652 9764 48692 23575
rect 49036 18752 49076 18761
rect 49036 16820 49076 18712
rect 50379 18332 50421 18341
rect 50379 18292 50380 18332
rect 50420 18292 50421 18332
rect 50379 18283 50421 18292
rect 50380 17249 50420 18283
rect 50379 17240 50421 17249
rect 50379 17200 50380 17240
rect 50420 17200 50421 17240
rect 50379 17191 50421 17200
rect 49036 16771 49076 16780
rect 50764 14804 50804 27364
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 51628 25220 51668 31396
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 54604 28580 54644 28589
rect 52108 28076 52148 28085
rect 51628 25171 51668 25180
rect 52012 27488 52052 27497
rect 51340 23960 51380 23969
rect 50859 23540 50901 23549
rect 50859 23500 50860 23540
rect 50900 23500 50901 23540
rect 50859 23491 50901 23500
rect 50764 14755 50804 14764
rect 49324 14636 49364 14645
rect 49324 13208 49364 14596
rect 49324 11024 49364 13168
rect 49324 10975 49364 10984
rect 48652 9715 48692 9724
rect 50860 8504 50900 23491
rect 51340 23120 51380 23920
rect 51723 23876 51765 23885
rect 51723 23836 51724 23876
rect 51764 23836 51765 23876
rect 51723 23827 51765 23836
rect 51724 23708 51764 23827
rect 51627 23456 51669 23465
rect 51627 23416 51628 23456
rect 51668 23416 51669 23456
rect 51627 23407 51669 23416
rect 51531 23204 51573 23213
rect 51531 23164 51532 23204
rect 51572 23164 51573 23204
rect 51531 23155 51573 23164
rect 51340 23071 51380 23080
rect 51339 18500 51381 18509
rect 51339 18460 51340 18500
rect 51380 18460 51381 18500
rect 51339 18451 51381 18460
rect 51340 18416 51380 18451
rect 51340 18365 51380 18376
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 51532 12368 51572 23155
rect 51628 21272 51668 23407
rect 51628 21223 51668 21232
rect 51532 12319 51572 12328
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 50860 8455 50900 8464
rect 48844 8336 48884 8345
rect 48844 7664 48884 8296
rect 48844 7615 48884 7624
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 48172 6187 48212 6196
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 51724 2624 51764 23668
rect 51819 23372 51861 23381
rect 51819 23332 51820 23372
rect 51860 23332 51861 23372
rect 51819 23323 51861 23332
rect 51820 22616 51860 23323
rect 51820 22567 51860 22576
rect 51916 18584 51956 18593
rect 51820 18500 51860 18509
rect 51820 16241 51860 18460
rect 51916 16829 51956 18544
rect 51915 16820 51957 16829
rect 51915 16780 51916 16820
rect 51956 16780 51957 16820
rect 51915 16771 51957 16780
rect 52012 16325 52052 27448
rect 52011 16316 52053 16325
rect 52011 16276 52012 16316
rect 52052 16276 52053 16316
rect 52011 16267 52053 16276
rect 51819 16232 51861 16241
rect 51819 16192 51820 16232
rect 51860 16192 51861 16232
rect 51819 16183 51861 16192
rect 51916 15980 51956 15989
rect 51916 13889 51956 15940
rect 52108 14813 52148 28036
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 52780 27992 52820 28001
rect 52780 27488 52820 27952
rect 52780 27439 52820 27448
rect 52972 27152 53012 27161
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 52875 26480 52917 26489
rect 52875 26440 52876 26480
rect 52916 26440 52917 26480
rect 52875 26431 52917 26440
rect 52204 26144 52244 26153
rect 52107 14804 52149 14813
rect 52107 14764 52108 14804
rect 52148 14764 52149 14804
rect 52107 14755 52149 14764
rect 51915 13880 51957 13889
rect 51915 13840 51916 13880
rect 51956 13840 51957 13880
rect 51915 13831 51957 13840
rect 51916 12872 51956 13831
rect 51916 12823 51956 12832
rect 52204 11948 52244 26104
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 52492 23288 52532 23297
rect 52492 22877 52532 23248
rect 52587 23120 52629 23129
rect 52587 23080 52588 23120
rect 52628 23080 52629 23120
rect 52587 23071 52629 23080
rect 52491 22868 52533 22877
rect 52491 22828 52492 22868
rect 52532 22828 52533 22868
rect 52491 22819 52533 22828
rect 52300 22196 52340 22205
rect 52300 20936 52340 22156
rect 52300 20887 52340 20896
rect 52492 20264 52532 22819
rect 52588 21608 52628 23071
rect 52588 21559 52628 21568
rect 52492 20215 52532 20224
rect 52299 17576 52341 17585
rect 52299 17536 52300 17576
rect 52340 17536 52341 17576
rect 52299 17527 52341 17536
rect 52300 17165 52340 17527
rect 52299 17156 52341 17165
rect 52299 17116 52300 17156
rect 52340 17116 52341 17156
rect 52299 17107 52341 17116
rect 52779 17156 52821 17165
rect 52779 17116 52780 17156
rect 52820 17116 52821 17156
rect 52779 17107 52821 17116
rect 52300 17022 52340 17107
rect 52587 17072 52629 17081
rect 52587 17032 52588 17072
rect 52628 17032 52629 17072
rect 52587 17023 52629 17032
rect 52780 17072 52820 17107
rect 52588 16938 52628 17023
rect 52780 17021 52820 17032
rect 52780 16232 52820 16241
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 52780 14132 52820 16192
rect 52876 14981 52916 26431
rect 52875 14972 52917 14981
rect 52875 14932 52876 14972
rect 52916 14932 52917 14972
rect 52875 14923 52917 14932
rect 52780 14083 52820 14092
rect 52972 13049 53012 27112
rect 53068 26564 53108 26573
rect 53068 14897 53108 26524
rect 54507 26480 54549 26489
rect 54507 26440 54508 26480
rect 54548 26440 54549 26480
rect 54507 26431 54549 26440
rect 54508 26346 54548 26431
rect 54604 23885 54644 28540
rect 59404 28580 59444 38200
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 72460 37400 72500 37409
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 69100 36896 69140 36905
rect 69100 36476 69140 36856
rect 69100 36427 69140 36436
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 67564 36308 67604 36317
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 67564 33956 67604 36268
rect 67564 33907 67604 33916
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 70636 32612 70676 32621
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 64012 29168 64052 29177
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 59404 28531 59444 28540
rect 64012 28496 64052 29128
rect 60172 28328 60212 28337
rect 58252 27656 58292 27665
rect 56715 26228 56757 26237
rect 56715 26188 56716 26228
rect 56756 26188 56757 26228
rect 56715 26179 56757 26188
rect 56716 26069 56756 26179
rect 56715 26060 56757 26069
rect 56715 26020 56716 26060
rect 56756 26020 56757 26060
rect 56715 26011 56757 26020
rect 54603 23876 54645 23885
rect 54603 23836 54604 23876
rect 54644 23836 54645 23876
rect 54603 23827 54645 23836
rect 54796 23792 54836 23801
rect 54796 23633 54836 23752
rect 55852 23792 55892 23803
rect 55852 23717 55892 23752
rect 56812 23792 56852 23801
rect 55851 23708 55893 23717
rect 55851 23668 55852 23708
rect 55892 23668 55893 23708
rect 55851 23659 55893 23668
rect 54795 23624 54837 23633
rect 54795 23584 54796 23624
rect 54836 23584 54837 23624
rect 54795 23575 54837 23584
rect 54796 23456 54836 23575
rect 56139 23540 56181 23549
rect 56139 23500 56140 23540
rect 56180 23500 56181 23540
rect 56139 23491 56181 23500
rect 54796 23407 54836 23416
rect 55659 23204 55701 23213
rect 55659 23164 55660 23204
rect 55700 23164 55701 23204
rect 55659 23155 55701 23164
rect 54411 23120 54453 23129
rect 54411 23080 54412 23120
rect 54452 23080 54453 23120
rect 54411 23071 54453 23080
rect 54412 22784 54452 23071
rect 55660 23070 55700 23155
rect 56140 23036 56180 23491
rect 56812 23465 56852 23752
rect 57292 23792 57332 23801
rect 56811 23456 56853 23465
rect 56811 23416 56812 23456
rect 56852 23416 56853 23456
rect 56811 23407 56853 23416
rect 57292 23381 57332 23752
rect 58252 23624 58292 27616
rect 60172 27404 60212 28288
rect 60172 27355 60212 27364
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 58539 27068 58581 27077
rect 58539 27028 58540 27068
rect 58580 27028 58581 27068
rect 58539 27019 58581 27028
rect 58540 26934 58580 27019
rect 58348 26900 58388 26909
rect 58348 25985 58388 26860
rect 60364 26900 60404 26909
rect 60364 26237 60404 26860
rect 64012 26312 64052 28456
rect 65164 28496 65204 28505
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 65164 27320 65204 28456
rect 65164 27271 65204 27280
rect 67564 27572 67604 27581
rect 67564 27077 67604 27532
rect 67563 27068 67605 27077
rect 67563 27028 67564 27068
rect 67604 27028 67605 27068
rect 67563 27019 67605 27028
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 64012 26263 64052 26272
rect 60363 26228 60405 26237
rect 60363 26188 60364 26228
rect 60404 26188 60405 26228
rect 60363 26179 60405 26188
rect 59404 26144 59444 26153
rect 58347 25976 58389 25985
rect 58347 25936 58348 25976
rect 58388 25936 58389 25976
rect 58347 25927 58389 25936
rect 59404 25892 59444 26104
rect 59404 25843 59444 25852
rect 60364 26060 60404 26069
rect 60364 25136 60404 26020
rect 60555 26060 60597 26069
rect 60555 26020 60556 26060
rect 60596 26020 60597 26060
rect 60555 26011 60597 26020
rect 60556 25926 60596 26011
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 60364 25087 60404 25096
rect 63916 25640 63956 25649
rect 63916 25052 63956 25600
rect 63916 24716 63956 25012
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 63916 24667 63956 24676
rect 70636 23792 70676 32572
rect 71980 31436 72020 31445
rect 71116 31184 71156 31193
rect 71116 30008 71156 31144
rect 71980 30596 72020 31396
rect 71116 29959 71156 29968
rect 71308 30176 71348 30185
rect 71308 29756 71348 30136
rect 71308 29707 71348 29716
rect 71404 28832 71444 28841
rect 71404 27320 71444 28792
rect 71404 27271 71444 27280
rect 71692 28076 71732 28085
rect 70636 23743 70676 23752
rect 71692 23792 71732 28036
rect 71980 27488 72020 30556
rect 72460 30260 72500 37360
rect 76972 37400 77012 37409
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 76876 36224 76916 36233
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 76352 34040 76720 34049
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 76876 33788 76916 36184
rect 75112 33284 75480 33293
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75112 33235 75480 33244
rect 76352 32528 76720 32537
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76352 32479 76720 32488
rect 76876 32276 76916 33748
rect 75112 31772 75480 31781
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75112 31723 75480 31732
rect 76876 31184 76916 32236
rect 76876 31135 76916 31144
rect 76352 31016 76720 31025
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76352 30967 76720 30976
rect 72460 30211 72500 30220
rect 75112 30260 75480 30269
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75112 30211 75480 30220
rect 76108 30260 76148 30269
rect 75112 28748 75480 28757
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75112 28699 75480 28708
rect 71980 26564 72020 27448
rect 75112 27236 75480 27245
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75112 27187 75480 27196
rect 71980 26515 72020 26524
rect 75112 25724 75480 25733
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75112 25675 75480 25684
rect 71692 23743 71732 23752
rect 76108 23792 76148 30220
rect 76352 29504 76720 29513
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76352 29455 76720 29464
rect 76352 27992 76720 28001
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76352 27943 76720 27952
rect 76352 26480 76720 26489
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76352 26431 76720 26440
rect 76352 24968 76720 24977
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76352 24919 76720 24928
rect 76108 23743 76148 23752
rect 76972 23792 77012 37360
rect 77452 32192 77492 32201
rect 77260 31268 77300 31277
rect 77260 30596 77300 31228
rect 77260 30260 77300 30556
rect 77260 30211 77300 30220
rect 76972 23743 77012 23752
rect 77452 23792 77492 32152
rect 77836 28748 77876 28757
rect 77836 25892 77876 28708
rect 77836 25843 77876 25852
rect 77452 23743 77492 23752
rect 79083 23792 79125 23801
rect 79083 23752 79084 23792
rect 79124 23752 79125 23792
rect 79083 23743 79125 23752
rect 79084 23658 79124 23743
rect 58252 23575 58292 23584
rect 60556 23624 60596 23633
rect 57291 23372 57333 23381
rect 57291 23332 57292 23372
rect 57332 23332 57333 23372
rect 57291 23323 57333 23332
rect 57675 23372 57717 23381
rect 57675 23332 57676 23372
rect 57716 23332 57717 23372
rect 57675 23323 57717 23332
rect 56811 23288 56853 23297
rect 56811 23248 56812 23288
rect 56852 23248 56853 23288
rect 56811 23239 56853 23248
rect 56812 23154 56852 23239
rect 56140 22987 56180 22996
rect 54700 22877 54740 22962
rect 54699 22868 54741 22877
rect 54699 22828 54700 22868
rect 54740 22828 54741 22868
rect 54699 22819 54741 22828
rect 54412 22735 54452 22744
rect 57676 22784 57716 23323
rect 57676 22735 57716 22744
rect 60556 22784 60596 23584
rect 60556 22735 60596 22744
rect 54316 17240 54356 17249
rect 54316 16829 54356 17200
rect 55083 17240 55125 17249
rect 55083 17200 55084 17240
rect 55124 17200 55125 17240
rect 55083 17191 55125 17200
rect 58252 17240 58292 17249
rect 54700 17072 54740 17083
rect 54700 16997 54740 17032
rect 54699 16988 54741 16997
rect 54699 16948 54700 16988
rect 54740 16948 54741 16988
rect 54699 16939 54741 16948
rect 54315 16820 54357 16829
rect 54315 16780 54316 16820
rect 54356 16780 54357 16820
rect 54315 16771 54357 16780
rect 55084 16232 55124 17191
rect 57868 17156 57908 17165
rect 57868 16745 57908 17116
rect 58252 16913 58292 17200
rect 75724 17240 75764 17249
rect 58251 16904 58293 16913
rect 58251 16864 58252 16904
rect 58292 16864 58293 16904
rect 58251 16855 58293 16864
rect 57867 16736 57909 16745
rect 57867 16696 57868 16736
rect 57908 16696 57909 16736
rect 57867 16687 57909 16696
rect 61707 16316 61749 16325
rect 61707 16276 61708 16316
rect 61748 16276 61749 16316
rect 61707 16267 61749 16276
rect 55084 16183 55124 16192
rect 58540 16232 58580 16241
rect 53067 14888 53109 14897
rect 53067 14848 53068 14888
rect 53108 14848 53109 14888
rect 53067 14839 53109 14848
rect 58540 14561 58580 16192
rect 61708 16182 61748 16267
rect 64971 16232 65013 16241
rect 64971 16192 64972 16232
rect 65012 16192 65013 16232
rect 64971 16183 65013 16192
rect 70156 16232 70196 16241
rect 64972 16098 65012 16183
rect 68524 16064 68564 16073
rect 60652 15812 60692 15821
rect 58923 14804 58965 14813
rect 58923 14764 58924 14804
rect 58964 14764 58965 14804
rect 58923 14755 58965 14764
rect 58539 14552 58581 14561
rect 58539 14512 58540 14552
rect 58580 14512 58581 14552
rect 58539 14503 58581 14512
rect 57772 14048 57812 14057
rect 57772 13889 57812 14008
rect 57867 13964 57909 13973
rect 57867 13924 57868 13964
rect 57908 13924 57909 13964
rect 57867 13915 57909 13924
rect 57771 13880 57813 13889
rect 57771 13840 57772 13880
rect 57812 13840 57813 13880
rect 57771 13831 57813 13840
rect 57868 13049 57908 13915
rect 52971 13040 53013 13049
rect 52971 13000 52972 13040
rect 53012 13000 53013 13040
rect 52971 12991 53013 13000
rect 57867 13040 57909 13049
rect 57867 13000 57868 13040
rect 57908 13000 57909 13040
rect 57867 12991 57909 13000
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 52204 11899 52244 11908
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 58924 10268 58964 14755
rect 60652 11948 60692 15772
rect 62956 15392 62996 15401
rect 63340 15392 63380 15401
rect 62996 15352 63340 15392
rect 62956 15343 62996 15352
rect 63340 15343 63380 15352
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 60748 15056 60788 15065
rect 60748 14897 60788 15016
rect 61899 14972 61941 14981
rect 61899 14932 61900 14972
rect 61940 14932 61941 14972
rect 61899 14923 61941 14932
rect 60747 14888 60789 14897
rect 60747 14848 60748 14888
rect 60788 14848 60789 14888
rect 60747 14839 60789 14848
rect 61900 14888 61940 14923
rect 60748 14720 60788 14839
rect 61900 14837 61940 14848
rect 67179 14804 67221 14813
rect 67179 14764 67180 14804
rect 67220 14764 67221 14804
rect 67179 14755 67221 14764
rect 60748 14671 60788 14680
rect 67180 14670 67220 14755
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 63916 13964 63956 13973
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 63532 12536 63572 12545
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 60652 11899 60692 11908
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 63532 10436 63572 12496
rect 63916 12536 63956 13924
rect 68524 13796 68564 16024
rect 68524 13747 68564 13756
rect 69100 16064 69140 16073
rect 68908 13040 68948 13049
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 63916 12487 63956 12496
rect 68908 11696 68948 13000
rect 68908 11647 68948 11656
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 63532 10387 63572 10396
rect 58924 10219 58964 10228
rect 69100 10100 69140 16024
rect 69195 13964 69237 13973
rect 69195 13924 69196 13964
rect 69236 13924 69237 13964
rect 69195 13915 69237 13924
rect 69196 13880 69236 13915
rect 69196 13829 69236 13840
rect 69100 10051 69140 10060
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 66316 8000 66356 8009
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 66316 5480 66356 7960
rect 66316 5431 66356 5440
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 70156 4472 70196 16192
rect 75724 16232 75764 17200
rect 78891 17072 78933 17081
rect 78891 17032 78892 17072
rect 78932 17032 78933 17072
rect 78891 17023 78933 17032
rect 78892 16241 78932 17023
rect 75112 15140 75480 15149
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75112 15091 75480 15100
rect 75112 13628 75480 13637
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75112 13579 75480 13588
rect 74860 13460 74900 13469
rect 74860 13124 74900 13420
rect 70539 11612 70581 11621
rect 70539 11572 70540 11612
rect 70580 11572 70581 11612
rect 70539 11563 70581 11572
rect 70540 11478 70580 11563
rect 74860 11360 74900 13084
rect 75112 12116 75480 12125
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75112 12067 75480 12076
rect 74860 11311 74900 11320
rect 75112 10604 75480 10613
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75112 10555 75480 10564
rect 75112 9092 75480 9101
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75112 9043 75480 9052
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 70156 4423 70196 4432
rect 71308 5648 71348 5657
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 71308 3716 71348 5608
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 51724 2575 51764 2584
rect 71308 2540 71348 3676
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 75724 2624 75764 16192
rect 77644 16232 77684 16241
rect 77356 16064 77396 16073
rect 76352 14384 76720 14393
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76352 14335 76720 14344
rect 76204 13208 76244 13217
rect 76204 11621 76244 13168
rect 76352 12872 76720 12881
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76352 12823 76720 12832
rect 76203 11612 76245 11621
rect 76203 11572 76204 11612
rect 76244 11572 76245 11612
rect 76203 11563 76245 11572
rect 76395 11612 76437 11621
rect 76395 11572 76396 11612
rect 76436 11572 76437 11612
rect 76395 11563 76437 11572
rect 76396 11478 76436 11563
rect 76352 11360 76720 11369
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76352 11311 76720 11320
rect 76352 9848 76720 9857
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76352 9799 76720 9808
rect 76204 9596 76244 9605
rect 76204 8420 76244 9556
rect 76204 8371 76244 8380
rect 76352 8336 76720 8345
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76352 8287 76720 8296
rect 76204 7412 76244 7421
rect 76204 6824 76244 7372
rect 76204 6775 76244 6784
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 76204 4388 76244 4397
rect 76204 3464 76244 4348
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 76204 3415 76244 3424
rect 75724 2575 75764 2584
rect 77356 2624 77396 16024
rect 77644 7160 77684 16192
rect 78891 16232 78933 16241
rect 78891 16192 78892 16232
rect 78932 16192 78933 16232
rect 78891 16183 78933 16192
rect 78892 16098 78932 16183
rect 77644 7111 77684 7120
rect 77356 2575 77396 2584
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 71308 2288 71348 2500
rect 71308 2239 71348 2248
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 38860 25936 38900 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 11692 23164 11732 23204
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 40876 26020 40916 26060
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 43180 26104 43220 26144
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 48172 23668 48212 23708
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 35404 18292 35444 18332
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 25516 17536 25556 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 43084 18460 43124 18500
rect 32812 16948 32852 16988
rect 36652 16864 36692 16904
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 29644 16780 29684 16820
rect 39724 16696 39764 16736
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 32332 14512 32372 14552
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 48652 23584 48692 23624
rect 50380 18292 50420 18332
rect 50380 17200 50420 17240
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 50860 23500 50900 23540
rect 51724 23836 51764 23876
rect 51628 23416 51668 23456
rect 51532 23164 51572 23204
rect 51340 18460 51380 18500
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 51820 23332 51860 23372
rect 51916 16780 51956 16820
rect 52012 16276 52052 16316
rect 51820 16192 51860 16232
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 52876 26440 52916 26480
rect 52108 14764 52148 14804
rect 51916 13840 51956 13880
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 52588 23080 52628 23120
rect 52492 22828 52532 22868
rect 52300 17536 52340 17576
rect 52300 17116 52340 17156
rect 52780 17116 52820 17156
rect 52588 17032 52628 17072
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 52876 14932 52916 14972
rect 54508 26440 54548 26480
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 56716 26188 56756 26228
rect 56716 26020 56756 26060
rect 54604 23836 54644 23876
rect 55852 23668 55892 23708
rect 54796 23584 54836 23624
rect 56140 23500 56180 23540
rect 55660 23164 55700 23204
rect 54412 23080 54452 23120
rect 56812 23416 56852 23456
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 58540 27028 58580 27068
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 67564 27028 67604 27068
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 60364 26188 60404 26228
rect 58348 25936 58388 25976
rect 60556 26020 60596 26060
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 79084 23752 79124 23792
rect 57292 23332 57332 23372
rect 57676 23332 57716 23372
rect 56812 23248 56852 23288
rect 54700 22828 54740 22868
rect 55084 17200 55124 17240
rect 54700 16948 54740 16988
rect 54316 16780 54356 16820
rect 58252 16864 58292 16904
rect 57868 16696 57908 16736
rect 61708 16276 61748 16316
rect 53068 14848 53108 14888
rect 64972 16192 65012 16232
rect 58924 14764 58964 14804
rect 58540 14512 58580 14552
rect 57868 13924 57908 13964
rect 57772 13840 57812 13880
rect 52972 13000 53012 13040
rect 57868 13000 57908 13040
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 61900 14932 61940 14972
rect 60748 14848 60788 14888
rect 67180 14764 67220 14804
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 69196 13924 69236 13964
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 78892 17032 78932 17072
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 70540 11572 70580 11612
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 76204 11572 76244 11612
rect 76396 11572 76436 11612
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 78892 16192 78932 16232
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 16343 38576 16390 38618
rect 16514 38576 16558 38618
rect 16682 38576 16729 38618
rect 16343 38536 16352 38576
rect 16514 38536 16516 38576
rect 16556 38536 16558 38576
rect 16720 38536 16729 38576
rect 16343 38494 16390 38536
rect 16514 38494 16558 38536
rect 16682 38494 16729 38536
rect 28343 38576 28390 38618
rect 28514 38576 28558 38618
rect 28682 38576 28729 38618
rect 28343 38536 28352 38576
rect 28514 38536 28516 38576
rect 28556 38536 28558 38576
rect 28720 38536 28729 38576
rect 28343 38494 28390 38536
rect 28514 38494 28558 38536
rect 28682 38494 28729 38536
rect 40343 38576 40390 38618
rect 40514 38576 40558 38618
rect 40682 38576 40729 38618
rect 40343 38536 40352 38576
rect 40514 38536 40516 38576
rect 40556 38536 40558 38576
rect 40720 38536 40729 38576
rect 40343 38494 40390 38536
rect 40514 38494 40558 38536
rect 40682 38494 40729 38536
rect 52343 38576 52390 38618
rect 52514 38576 52558 38618
rect 52682 38576 52729 38618
rect 52343 38536 52352 38576
rect 52514 38536 52516 38576
rect 52556 38536 52558 38576
rect 52720 38536 52729 38576
rect 52343 38494 52390 38536
rect 52514 38494 52558 38536
rect 52682 38494 52729 38536
rect 64343 38576 64390 38618
rect 64514 38576 64558 38618
rect 64682 38576 64729 38618
rect 64343 38536 64352 38576
rect 64514 38536 64516 38576
rect 64556 38536 64558 38576
rect 64720 38536 64729 38576
rect 64343 38494 64390 38536
rect 64514 38494 64558 38536
rect 64682 38494 64729 38536
rect 76343 38576 76390 38618
rect 76514 38576 76558 38618
rect 76682 38576 76729 38618
rect 76343 38536 76352 38576
rect 76514 38536 76516 38576
rect 76556 38536 76558 38576
rect 76720 38536 76729 38576
rect 76343 38494 76390 38536
rect 76514 38494 76558 38536
rect 76682 38494 76729 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 15103 37820 15150 37862
rect 15274 37820 15318 37862
rect 15442 37820 15489 37862
rect 15103 37780 15112 37820
rect 15274 37780 15276 37820
rect 15316 37780 15318 37820
rect 15480 37780 15489 37820
rect 15103 37738 15150 37780
rect 15274 37738 15318 37780
rect 15442 37738 15489 37780
rect 27103 37820 27150 37862
rect 27274 37820 27318 37862
rect 27442 37820 27489 37862
rect 27103 37780 27112 37820
rect 27274 37780 27276 37820
rect 27316 37780 27318 37820
rect 27480 37780 27489 37820
rect 27103 37738 27150 37780
rect 27274 37738 27318 37780
rect 27442 37738 27489 37780
rect 39103 37820 39150 37862
rect 39274 37820 39318 37862
rect 39442 37820 39489 37862
rect 39103 37780 39112 37820
rect 39274 37780 39276 37820
rect 39316 37780 39318 37820
rect 39480 37780 39489 37820
rect 39103 37738 39150 37780
rect 39274 37738 39318 37780
rect 39442 37738 39489 37780
rect 51103 37820 51150 37862
rect 51274 37820 51318 37862
rect 51442 37820 51489 37862
rect 51103 37780 51112 37820
rect 51274 37780 51276 37820
rect 51316 37780 51318 37820
rect 51480 37780 51489 37820
rect 51103 37738 51150 37780
rect 51274 37738 51318 37780
rect 51442 37738 51489 37780
rect 63103 37820 63150 37862
rect 63274 37820 63318 37862
rect 63442 37820 63489 37862
rect 63103 37780 63112 37820
rect 63274 37780 63276 37820
rect 63316 37780 63318 37820
rect 63480 37780 63489 37820
rect 63103 37738 63150 37780
rect 63274 37738 63318 37780
rect 63442 37738 63489 37780
rect 75103 37820 75150 37862
rect 75274 37820 75318 37862
rect 75442 37820 75489 37862
rect 75103 37780 75112 37820
rect 75274 37780 75276 37820
rect 75316 37780 75318 37820
rect 75480 37780 75489 37820
rect 75103 37738 75150 37780
rect 75274 37738 75318 37780
rect 75442 37738 75489 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 16343 37064 16390 37106
rect 16514 37064 16558 37106
rect 16682 37064 16729 37106
rect 16343 37024 16352 37064
rect 16514 37024 16516 37064
rect 16556 37024 16558 37064
rect 16720 37024 16729 37064
rect 16343 36982 16390 37024
rect 16514 36982 16558 37024
rect 16682 36982 16729 37024
rect 28343 37064 28390 37106
rect 28514 37064 28558 37106
rect 28682 37064 28729 37106
rect 28343 37024 28352 37064
rect 28514 37024 28516 37064
rect 28556 37024 28558 37064
rect 28720 37024 28729 37064
rect 28343 36982 28390 37024
rect 28514 36982 28558 37024
rect 28682 36982 28729 37024
rect 40343 37064 40390 37106
rect 40514 37064 40558 37106
rect 40682 37064 40729 37106
rect 40343 37024 40352 37064
rect 40514 37024 40516 37064
rect 40556 37024 40558 37064
rect 40720 37024 40729 37064
rect 40343 36982 40390 37024
rect 40514 36982 40558 37024
rect 40682 36982 40729 37024
rect 52343 37064 52390 37106
rect 52514 37064 52558 37106
rect 52682 37064 52729 37106
rect 52343 37024 52352 37064
rect 52514 37024 52516 37064
rect 52556 37024 52558 37064
rect 52720 37024 52729 37064
rect 52343 36982 52390 37024
rect 52514 36982 52558 37024
rect 52682 36982 52729 37024
rect 64343 37064 64390 37106
rect 64514 37064 64558 37106
rect 64682 37064 64729 37106
rect 64343 37024 64352 37064
rect 64514 37024 64516 37064
rect 64556 37024 64558 37064
rect 64720 37024 64729 37064
rect 64343 36982 64390 37024
rect 64514 36982 64558 37024
rect 64682 36982 64729 37024
rect 76343 37064 76390 37106
rect 76514 37064 76558 37106
rect 76682 37064 76729 37106
rect 76343 37024 76352 37064
rect 76514 37024 76516 37064
rect 76556 37024 76558 37064
rect 76720 37024 76729 37064
rect 76343 36982 76390 37024
rect 76514 36982 76558 37024
rect 76682 36982 76729 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 15103 36308 15150 36350
rect 15274 36308 15318 36350
rect 15442 36308 15489 36350
rect 15103 36268 15112 36308
rect 15274 36268 15276 36308
rect 15316 36268 15318 36308
rect 15480 36268 15489 36308
rect 15103 36226 15150 36268
rect 15274 36226 15318 36268
rect 15442 36226 15489 36268
rect 27103 36308 27150 36350
rect 27274 36308 27318 36350
rect 27442 36308 27489 36350
rect 27103 36268 27112 36308
rect 27274 36268 27276 36308
rect 27316 36268 27318 36308
rect 27480 36268 27489 36308
rect 27103 36226 27150 36268
rect 27274 36226 27318 36268
rect 27442 36226 27489 36268
rect 39103 36308 39150 36350
rect 39274 36308 39318 36350
rect 39442 36308 39489 36350
rect 39103 36268 39112 36308
rect 39274 36268 39276 36308
rect 39316 36268 39318 36308
rect 39480 36268 39489 36308
rect 39103 36226 39150 36268
rect 39274 36226 39318 36268
rect 39442 36226 39489 36268
rect 51103 36308 51150 36350
rect 51274 36308 51318 36350
rect 51442 36308 51489 36350
rect 51103 36268 51112 36308
rect 51274 36268 51276 36308
rect 51316 36268 51318 36308
rect 51480 36268 51489 36308
rect 51103 36226 51150 36268
rect 51274 36226 51318 36268
rect 51442 36226 51489 36268
rect 63103 36308 63150 36350
rect 63274 36308 63318 36350
rect 63442 36308 63489 36350
rect 63103 36268 63112 36308
rect 63274 36268 63276 36308
rect 63316 36268 63318 36308
rect 63480 36268 63489 36308
rect 63103 36226 63150 36268
rect 63274 36226 63318 36268
rect 63442 36226 63489 36268
rect 75103 36308 75150 36350
rect 75274 36308 75318 36350
rect 75442 36308 75489 36350
rect 75103 36268 75112 36308
rect 75274 36268 75276 36308
rect 75316 36268 75318 36308
rect 75480 36268 75489 36308
rect 75103 36226 75150 36268
rect 75274 36226 75318 36268
rect 75442 36226 75489 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 16343 35552 16390 35594
rect 16514 35552 16558 35594
rect 16682 35552 16729 35594
rect 16343 35512 16352 35552
rect 16514 35512 16516 35552
rect 16556 35512 16558 35552
rect 16720 35512 16729 35552
rect 16343 35470 16390 35512
rect 16514 35470 16558 35512
rect 16682 35470 16729 35512
rect 28343 35552 28390 35594
rect 28514 35552 28558 35594
rect 28682 35552 28729 35594
rect 28343 35512 28352 35552
rect 28514 35512 28516 35552
rect 28556 35512 28558 35552
rect 28720 35512 28729 35552
rect 28343 35470 28390 35512
rect 28514 35470 28558 35512
rect 28682 35470 28729 35512
rect 40343 35552 40390 35594
rect 40514 35552 40558 35594
rect 40682 35552 40729 35594
rect 40343 35512 40352 35552
rect 40514 35512 40516 35552
rect 40556 35512 40558 35552
rect 40720 35512 40729 35552
rect 40343 35470 40390 35512
rect 40514 35470 40558 35512
rect 40682 35470 40729 35512
rect 52343 35552 52390 35594
rect 52514 35552 52558 35594
rect 52682 35552 52729 35594
rect 52343 35512 52352 35552
rect 52514 35512 52516 35552
rect 52556 35512 52558 35552
rect 52720 35512 52729 35552
rect 52343 35470 52390 35512
rect 52514 35470 52558 35512
rect 52682 35470 52729 35512
rect 64343 35552 64390 35594
rect 64514 35552 64558 35594
rect 64682 35552 64729 35594
rect 64343 35512 64352 35552
rect 64514 35512 64516 35552
rect 64556 35512 64558 35552
rect 64720 35512 64729 35552
rect 64343 35470 64390 35512
rect 64514 35470 64558 35512
rect 64682 35470 64729 35512
rect 76343 35552 76390 35594
rect 76514 35552 76558 35594
rect 76682 35552 76729 35594
rect 76343 35512 76352 35552
rect 76514 35512 76516 35552
rect 76556 35512 76558 35552
rect 76720 35512 76729 35552
rect 76343 35470 76390 35512
rect 76514 35470 76558 35512
rect 76682 35470 76729 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 15103 34796 15150 34838
rect 15274 34796 15318 34838
rect 15442 34796 15489 34838
rect 15103 34756 15112 34796
rect 15274 34756 15276 34796
rect 15316 34756 15318 34796
rect 15480 34756 15489 34796
rect 15103 34714 15150 34756
rect 15274 34714 15318 34756
rect 15442 34714 15489 34756
rect 27103 34796 27150 34838
rect 27274 34796 27318 34838
rect 27442 34796 27489 34838
rect 27103 34756 27112 34796
rect 27274 34756 27276 34796
rect 27316 34756 27318 34796
rect 27480 34756 27489 34796
rect 27103 34714 27150 34756
rect 27274 34714 27318 34756
rect 27442 34714 27489 34756
rect 39103 34796 39150 34838
rect 39274 34796 39318 34838
rect 39442 34796 39489 34838
rect 39103 34756 39112 34796
rect 39274 34756 39276 34796
rect 39316 34756 39318 34796
rect 39480 34756 39489 34796
rect 39103 34714 39150 34756
rect 39274 34714 39318 34756
rect 39442 34714 39489 34756
rect 51103 34796 51150 34838
rect 51274 34796 51318 34838
rect 51442 34796 51489 34838
rect 51103 34756 51112 34796
rect 51274 34756 51276 34796
rect 51316 34756 51318 34796
rect 51480 34756 51489 34796
rect 51103 34714 51150 34756
rect 51274 34714 51318 34756
rect 51442 34714 51489 34756
rect 63103 34796 63150 34838
rect 63274 34796 63318 34838
rect 63442 34796 63489 34838
rect 63103 34756 63112 34796
rect 63274 34756 63276 34796
rect 63316 34756 63318 34796
rect 63480 34756 63489 34796
rect 63103 34714 63150 34756
rect 63274 34714 63318 34756
rect 63442 34714 63489 34756
rect 75103 34796 75150 34838
rect 75274 34796 75318 34838
rect 75442 34796 75489 34838
rect 75103 34756 75112 34796
rect 75274 34756 75276 34796
rect 75316 34756 75318 34796
rect 75480 34756 75489 34796
rect 75103 34714 75150 34756
rect 75274 34714 75318 34756
rect 75442 34714 75489 34756
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 16343 34040 16390 34082
rect 16514 34040 16558 34082
rect 16682 34040 16729 34082
rect 16343 34000 16352 34040
rect 16514 34000 16516 34040
rect 16556 34000 16558 34040
rect 16720 34000 16729 34040
rect 16343 33958 16390 34000
rect 16514 33958 16558 34000
rect 16682 33958 16729 34000
rect 28343 34040 28390 34082
rect 28514 34040 28558 34082
rect 28682 34040 28729 34082
rect 28343 34000 28352 34040
rect 28514 34000 28516 34040
rect 28556 34000 28558 34040
rect 28720 34000 28729 34040
rect 28343 33958 28390 34000
rect 28514 33958 28558 34000
rect 28682 33958 28729 34000
rect 40343 34040 40390 34082
rect 40514 34040 40558 34082
rect 40682 34040 40729 34082
rect 40343 34000 40352 34040
rect 40514 34000 40516 34040
rect 40556 34000 40558 34040
rect 40720 34000 40729 34040
rect 40343 33958 40390 34000
rect 40514 33958 40558 34000
rect 40682 33958 40729 34000
rect 52343 34040 52390 34082
rect 52514 34040 52558 34082
rect 52682 34040 52729 34082
rect 52343 34000 52352 34040
rect 52514 34000 52516 34040
rect 52556 34000 52558 34040
rect 52720 34000 52729 34040
rect 52343 33958 52390 34000
rect 52514 33958 52558 34000
rect 52682 33958 52729 34000
rect 64343 34040 64390 34082
rect 64514 34040 64558 34082
rect 64682 34040 64729 34082
rect 64343 34000 64352 34040
rect 64514 34000 64516 34040
rect 64556 34000 64558 34040
rect 64720 34000 64729 34040
rect 64343 33958 64390 34000
rect 64514 33958 64558 34000
rect 64682 33958 64729 34000
rect 76343 34040 76390 34082
rect 76514 34040 76558 34082
rect 76682 34040 76729 34082
rect 76343 34000 76352 34040
rect 76514 34000 76516 34040
rect 76556 34000 76558 34040
rect 76720 34000 76729 34040
rect 76343 33958 76390 34000
rect 76514 33958 76558 34000
rect 76682 33958 76729 34000
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 15103 33284 15150 33326
rect 15274 33284 15318 33326
rect 15442 33284 15489 33326
rect 15103 33244 15112 33284
rect 15274 33244 15276 33284
rect 15316 33244 15318 33284
rect 15480 33244 15489 33284
rect 15103 33202 15150 33244
rect 15274 33202 15318 33244
rect 15442 33202 15489 33244
rect 27103 33284 27150 33326
rect 27274 33284 27318 33326
rect 27442 33284 27489 33326
rect 27103 33244 27112 33284
rect 27274 33244 27276 33284
rect 27316 33244 27318 33284
rect 27480 33244 27489 33284
rect 27103 33202 27150 33244
rect 27274 33202 27318 33244
rect 27442 33202 27489 33244
rect 39103 33284 39150 33326
rect 39274 33284 39318 33326
rect 39442 33284 39489 33326
rect 39103 33244 39112 33284
rect 39274 33244 39276 33284
rect 39316 33244 39318 33284
rect 39480 33244 39489 33284
rect 39103 33202 39150 33244
rect 39274 33202 39318 33244
rect 39442 33202 39489 33244
rect 51103 33284 51150 33326
rect 51274 33284 51318 33326
rect 51442 33284 51489 33326
rect 51103 33244 51112 33284
rect 51274 33244 51276 33284
rect 51316 33244 51318 33284
rect 51480 33244 51489 33284
rect 51103 33202 51150 33244
rect 51274 33202 51318 33244
rect 51442 33202 51489 33244
rect 63103 33284 63150 33326
rect 63274 33284 63318 33326
rect 63442 33284 63489 33326
rect 63103 33244 63112 33284
rect 63274 33244 63276 33284
rect 63316 33244 63318 33284
rect 63480 33244 63489 33284
rect 63103 33202 63150 33244
rect 63274 33202 63318 33244
rect 63442 33202 63489 33244
rect 75103 33284 75150 33326
rect 75274 33284 75318 33326
rect 75442 33284 75489 33326
rect 75103 33244 75112 33284
rect 75274 33244 75276 33284
rect 75316 33244 75318 33284
rect 75480 33244 75489 33284
rect 75103 33202 75150 33244
rect 75274 33202 75318 33244
rect 75442 33202 75489 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 16343 32528 16390 32570
rect 16514 32528 16558 32570
rect 16682 32528 16729 32570
rect 16343 32488 16352 32528
rect 16514 32488 16516 32528
rect 16556 32488 16558 32528
rect 16720 32488 16729 32528
rect 16343 32446 16390 32488
rect 16514 32446 16558 32488
rect 16682 32446 16729 32488
rect 28343 32528 28390 32570
rect 28514 32528 28558 32570
rect 28682 32528 28729 32570
rect 28343 32488 28352 32528
rect 28514 32488 28516 32528
rect 28556 32488 28558 32528
rect 28720 32488 28729 32528
rect 28343 32446 28390 32488
rect 28514 32446 28558 32488
rect 28682 32446 28729 32488
rect 40343 32528 40390 32570
rect 40514 32528 40558 32570
rect 40682 32528 40729 32570
rect 40343 32488 40352 32528
rect 40514 32488 40516 32528
rect 40556 32488 40558 32528
rect 40720 32488 40729 32528
rect 40343 32446 40390 32488
rect 40514 32446 40558 32488
rect 40682 32446 40729 32488
rect 52343 32528 52390 32570
rect 52514 32528 52558 32570
rect 52682 32528 52729 32570
rect 52343 32488 52352 32528
rect 52514 32488 52516 32528
rect 52556 32488 52558 32528
rect 52720 32488 52729 32528
rect 52343 32446 52390 32488
rect 52514 32446 52558 32488
rect 52682 32446 52729 32488
rect 64343 32528 64390 32570
rect 64514 32528 64558 32570
rect 64682 32528 64729 32570
rect 64343 32488 64352 32528
rect 64514 32488 64516 32528
rect 64556 32488 64558 32528
rect 64720 32488 64729 32528
rect 64343 32446 64390 32488
rect 64514 32446 64558 32488
rect 64682 32446 64729 32488
rect 76343 32528 76390 32570
rect 76514 32528 76558 32570
rect 76682 32528 76729 32570
rect 76343 32488 76352 32528
rect 76514 32488 76516 32528
rect 76556 32488 76558 32528
rect 76720 32488 76729 32528
rect 76343 32446 76390 32488
rect 76514 32446 76558 32488
rect 76682 32446 76729 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 15103 31772 15150 31814
rect 15274 31772 15318 31814
rect 15442 31772 15489 31814
rect 15103 31732 15112 31772
rect 15274 31732 15276 31772
rect 15316 31732 15318 31772
rect 15480 31732 15489 31772
rect 15103 31690 15150 31732
rect 15274 31690 15318 31732
rect 15442 31690 15489 31732
rect 27103 31772 27150 31814
rect 27274 31772 27318 31814
rect 27442 31772 27489 31814
rect 27103 31732 27112 31772
rect 27274 31732 27276 31772
rect 27316 31732 27318 31772
rect 27480 31732 27489 31772
rect 27103 31690 27150 31732
rect 27274 31690 27318 31732
rect 27442 31690 27489 31732
rect 39103 31772 39150 31814
rect 39274 31772 39318 31814
rect 39442 31772 39489 31814
rect 39103 31732 39112 31772
rect 39274 31732 39276 31772
rect 39316 31732 39318 31772
rect 39480 31732 39489 31772
rect 39103 31690 39150 31732
rect 39274 31690 39318 31732
rect 39442 31690 39489 31732
rect 51103 31772 51150 31814
rect 51274 31772 51318 31814
rect 51442 31772 51489 31814
rect 51103 31732 51112 31772
rect 51274 31732 51276 31772
rect 51316 31732 51318 31772
rect 51480 31732 51489 31772
rect 51103 31690 51150 31732
rect 51274 31690 51318 31732
rect 51442 31690 51489 31732
rect 63103 31772 63150 31814
rect 63274 31772 63318 31814
rect 63442 31772 63489 31814
rect 63103 31732 63112 31772
rect 63274 31732 63276 31772
rect 63316 31732 63318 31772
rect 63480 31732 63489 31772
rect 63103 31690 63150 31732
rect 63274 31690 63318 31732
rect 63442 31690 63489 31732
rect 75103 31772 75150 31814
rect 75274 31772 75318 31814
rect 75442 31772 75489 31814
rect 75103 31732 75112 31772
rect 75274 31732 75276 31772
rect 75316 31732 75318 31772
rect 75480 31732 75489 31772
rect 75103 31690 75150 31732
rect 75274 31690 75318 31732
rect 75442 31690 75489 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 16343 31016 16390 31058
rect 16514 31016 16558 31058
rect 16682 31016 16729 31058
rect 16343 30976 16352 31016
rect 16514 30976 16516 31016
rect 16556 30976 16558 31016
rect 16720 30976 16729 31016
rect 16343 30934 16390 30976
rect 16514 30934 16558 30976
rect 16682 30934 16729 30976
rect 28343 31016 28390 31058
rect 28514 31016 28558 31058
rect 28682 31016 28729 31058
rect 28343 30976 28352 31016
rect 28514 30976 28516 31016
rect 28556 30976 28558 31016
rect 28720 30976 28729 31016
rect 28343 30934 28390 30976
rect 28514 30934 28558 30976
rect 28682 30934 28729 30976
rect 40343 31016 40390 31058
rect 40514 31016 40558 31058
rect 40682 31016 40729 31058
rect 40343 30976 40352 31016
rect 40514 30976 40516 31016
rect 40556 30976 40558 31016
rect 40720 30976 40729 31016
rect 40343 30934 40390 30976
rect 40514 30934 40558 30976
rect 40682 30934 40729 30976
rect 52343 31016 52390 31058
rect 52514 31016 52558 31058
rect 52682 31016 52729 31058
rect 52343 30976 52352 31016
rect 52514 30976 52516 31016
rect 52556 30976 52558 31016
rect 52720 30976 52729 31016
rect 52343 30934 52390 30976
rect 52514 30934 52558 30976
rect 52682 30934 52729 30976
rect 64343 31016 64390 31058
rect 64514 31016 64558 31058
rect 64682 31016 64729 31058
rect 64343 30976 64352 31016
rect 64514 30976 64516 31016
rect 64556 30976 64558 31016
rect 64720 30976 64729 31016
rect 64343 30934 64390 30976
rect 64514 30934 64558 30976
rect 64682 30934 64729 30976
rect 76343 31016 76390 31058
rect 76514 31016 76558 31058
rect 76682 31016 76729 31058
rect 76343 30976 76352 31016
rect 76514 30976 76516 31016
rect 76556 30976 76558 31016
rect 76720 30976 76729 31016
rect 76343 30934 76390 30976
rect 76514 30934 76558 30976
rect 76682 30934 76729 30976
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 15103 30260 15150 30302
rect 15274 30260 15318 30302
rect 15442 30260 15489 30302
rect 15103 30220 15112 30260
rect 15274 30220 15276 30260
rect 15316 30220 15318 30260
rect 15480 30220 15489 30260
rect 15103 30178 15150 30220
rect 15274 30178 15318 30220
rect 15442 30178 15489 30220
rect 27103 30260 27150 30302
rect 27274 30260 27318 30302
rect 27442 30260 27489 30302
rect 27103 30220 27112 30260
rect 27274 30220 27276 30260
rect 27316 30220 27318 30260
rect 27480 30220 27489 30260
rect 27103 30178 27150 30220
rect 27274 30178 27318 30220
rect 27442 30178 27489 30220
rect 39103 30260 39150 30302
rect 39274 30260 39318 30302
rect 39442 30260 39489 30302
rect 39103 30220 39112 30260
rect 39274 30220 39276 30260
rect 39316 30220 39318 30260
rect 39480 30220 39489 30260
rect 39103 30178 39150 30220
rect 39274 30178 39318 30220
rect 39442 30178 39489 30220
rect 51103 30260 51150 30302
rect 51274 30260 51318 30302
rect 51442 30260 51489 30302
rect 51103 30220 51112 30260
rect 51274 30220 51276 30260
rect 51316 30220 51318 30260
rect 51480 30220 51489 30260
rect 51103 30178 51150 30220
rect 51274 30178 51318 30220
rect 51442 30178 51489 30220
rect 63103 30260 63150 30302
rect 63274 30260 63318 30302
rect 63442 30260 63489 30302
rect 63103 30220 63112 30260
rect 63274 30220 63276 30260
rect 63316 30220 63318 30260
rect 63480 30220 63489 30260
rect 63103 30178 63150 30220
rect 63274 30178 63318 30220
rect 63442 30178 63489 30220
rect 75103 30260 75150 30302
rect 75274 30260 75318 30302
rect 75442 30260 75489 30302
rect 75103 30220 75112 30260
rect 75274 30220 75276 30260
rect 75316 30220 75318 30260
rect 75480 30220 75489 30260
rect 75103 30178 75150 30220
rect 75274 30178 75318 30220
rect 75442 30178 75489 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 16343 29504 16390 29546
rect 16514 29504 16558 29546
rect 16682 29504 16729 29546
rect 16343 29464 16352 29504
rect 16514 29464 16516 29504
rect 16556 29464 16558 29504
rect 16720 29464 16729 29504
rect 16343 29422 16390 29464
rect 16514 29422 16558 29464
rect 16682 29422 16729 29464
rect 28343 29504 28390 29546
rect 28514 29504 28558 29546
rect 28682 29504 28729 29546
rect 28343 29464 28352 29504
rect 28514 29464 28516 29504
rect 28556 29464 28558 29504
rect 28720 29464 28729 29504
rect 28343 29422 28390 29464
rect 28514 29422 28558 29464
rect 28682 29422 28729 29464
rect 40343 29504 40390 29546
rect 40514 29504 40558 29546
rect 40682 29504 40729 29546
rect 40343 29464 40352 29504
rect 40514 29464 40516 29504
rect 40556 29464 40558 29504
rect 40720 29464 40729 29504
rect 40343 29422 40390 29464
rect 40514 29422 40558 29464
rect 40682 29422 40729 29464
rect 52343 29504 52390 29546
rect 52514 29504 52558 29546
rect 52682 29504 52729 29546
rect 52343 29464 52352 29504
rect 52514 29464 52516 29504
rect 52556 29464 52558 29504
rect 52720 29464 52729 29504
rect 52343 29422 52390 29464
rect 52514 29422 52558 29464
rect 52682 29422 52729 29464
rect 64343 29504 64390 29546
rect 64514 29504 64558 29546
rect 64682 29504 64729 29546
rect 64343 29464 64352 29504
rect 64514 29464 64516 29504
rect 64556 29464 64558 29504
rect 64720 29464 64729 29504
rect 64343 29422 64390 29464
rect 64514 29422 64558 29464
rect 64682 29422 64729 29464
rect 76343 29504 76390 29546
rect 76514 29504 76558 29546
rect 76682 29504 76729 29546
rect 76343 29464 76352 29504
rect 76514 29464 76516 29504
rect 76556 29464 76558 29504
rect 76720 29464 76729 29504
rect 76343 29422 76390 29464
rect 76514 29422 76558 29464
rect 76682 29422 76729 29464
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 15103 28748 15150 28790
rect 15274 28748 15318 28790
rect 15442 28748 15489 28790
rect 15103 28708 15112 28748
rect 15274 28708 15276 28748
rect 15316 28708 15318 28748
rect 15480 28708 15489 28748
rect 15103 28666 15150 28708
rect 15274 28666 15318 28708
rect 15442 28666 15489 28708
rect 27103 28748 27150 28790
rect 27274 28748 27318 28790
rect 27442 28748 27489 28790
rect 27103 28708 27112 28748
rect 27274 28708 27276 28748
rect 27316 28708 27318 28748
rect 27480 28708 27489 28748
rect 27103 28666 27150 28708
rect 27274 28666 27318 28708
rect 27442 28666 27489 28708
rect 39103 28748 39150 28790
rect 39274 28748 39318 28790
rect 39442 28748 39489 28790
rect 39103 28708 39112 28748
rect 39274 28708 39276 28748
rect 39316 28708 39318 28748
rect 39480 28708 39489 28748
rect 39103 28666 39150 28708
rect 39274 28666 39318 28708
rect 39442 28666 39489 28708
rect 51103 28748 51150 28790
rect 51274 28748 51318 28790
rect 51442 28748 51489 28790
rect 51103 28708 51112 28748
rect 51274 28708 51276 28748
rect 51316 28708 51318 28748
rect 51480 28708 51489 28748
rect 51103 28666 51150 28708
rect 51274 28666 51318 28708
rect 51442 28666 51489 28708
rect 63103 28748 63150 28790
rect 63274 28748 63318 28790
rect 63442 28748 63489 28790
rect 63103 28708 63112 28748
rect 63274 28708 63276 28748
rect 63316 28708 63318 28748
rect 63480 28708 63489 28748
rect 63103 28666 63150 28708
rect 63274 28666 63318 28708
rect 63442 28666 63489 28708
rect 75103 28748 75150 28790
rect 75274 28748 75318 28790
rect 75442 28748 75489 28790
rect 75103 28708 75112 28748
rect 75274 28708 75276 28748
rect 75316 28708 75318 28748
rect 75480 28708 75489 28748
rect 75103 28666 75150 28708
rect 75274 28666 75318 28708
rect 75442 28666 75489 28708
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 16343 27992 16390 28034
rect 16514 27992 16558 28034
rect 16682 27992 16729 28034
rect 16343 27952 16352 27992
rect 16514 27952 16516 27992
rect 16556 27952 16558 27992
rect 16720 27952 16729 27992
rect 16343 27910 16390 27952
rect 16514 27910 16558 27952
rect 16682 27910 16729 27952
rect 28343 27992 28390 28034
rect 28514 27992 28558 28034
rect 28682 27992 28729 28034
rect 28343 27952 28352 27992
rect 28514 27952 28516 27992
rect 28556 27952 28558 27992
rect 28720 27952 28729 27992
rect 28343 27910 28390 27952
rect 28514 27910 28558 27952
rect 28682 27910 28729 27952
rect 40343 27992 40390 28034
rect 40514 27992 40558 28034
rect 40682 27992 40729 28034
rect 40343 27952 40352 27992
rect 40514 27952 40516 27992
rect 40556 27952 40558 27992
rect 40720 27952 40729 27992
rect 40343 27910 40390 27952
rect 40514 27910 40558 27952
rect 40682 27910 40729 27952
rect 52343 27992 52390 28034
rect 52514 27992 52558 28034
rect 52682 27992 52729 28034
rect 52343 27952 52352 27992
rect 52514 27952 52516 27992
rect 52556 27952 52558 27992
rect 52720 27952 52729 27992
rect 52343 27910 52390 27952
rect 52514 27910 52558 27952
rect 52682 27910 52729 27952
rect 64343 27992 64390 28034
rect 64514 27992 64558 28034
rect 64682 27992 64729 28034
rect 64343 27952 64352 27992
rect 64514 27952 64516 27992
rect 64556 27952 64558 27992
rect 64720 27952 64729 27992
rect 64343 27910 64390 27952
rect 64514 27910 64558 27952
rect 64682 27910 64729 27952
rect 76343 27992 76390 28034
rect 76514 27992 76558 28034
rect 76682 27992 76729 28034
rect 76343 27952 76352 27992
rect 76514 27952 76516 27992
rect 76556 27952 76558 27992
rect 76720 27952 76729 27992
rect 76343 27910 76390 27952
rect 76514 27910 76558 27952
rect 76682 27910 76729 27952
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 15103 27236 15150 27278
rect 15274 27236 15318 27278
rect 15442 27236 15489 27278
rect 15103 27196 15112 27236
rect 15274 27196 15276 27236
rect 15316 27196 15318 27236
rect 15480 27196 15489 27236
rect 15103 27154 15150 27196
rect 15274 27154 15318 27196
rect 15442 27154 15489 27196
rect 27103 27236 27150 27278
rect 27274 27236 27318 27278
rect 27442 27236 27489 27278
rect 27103 27196 27112 27236
rect 27274 27196 27276 27236
rect 27316 27196 27318 27236
rect 27480 27196 27489 27236
rect 27103 27154 27150 27196
rect 27274 27154 27318 27196
rect 27442 27154 27489 27196
rect 39103 27236 39150 27278
rect 39274 27236 39318 27278
rect 39442 27236 39489 27278
rect 39103 27196 39112 27236
rect 39274 27196 39276 27236
rect 39316 27196 39318 27236
rect 39480 27196 39489 27236
rect 39103 27154 39150 27196
rect 39274 27154 39318 27196
rect 39442 27154 39489 27196
rect 51103 27236 51150 27278
rect 51274 27236 51318 27278
rect 51442 27236 51489 27278
rect 51103 27196 51112 27236
rect 51274 27196 51276 27236
rect 51316 27196 51318 27236
rect 51480 27196 51489 27236
rect 51103 27154 51150 27196
rect 51274 27154 51318 27196
rect 51442 27154 51489 27196
rect 63103 27236 63150 27278
rect 63274 27236 63318 27278
rect 63442 27236 63489 27278
rect 63103 27196 63112 27236
rect 63274 27196 63276 27236
rect 63316 27196 63318 27236
rect 63480 27196 63489 27236
rect 63103 27154 63150 27196
rect 63274 27154 63318 27196
rect 63442 27154 63489 27196
rect 75103 27236 75150 27278
rect 75274 27236 75318 27278
rect 75442 27236 75489 27278
rect 75103 27196 75112 27236
rect 75274 27196 75276 27236
rect 75316 27196 75318 27236
rect 75480 27196 75489 27236
rect 75103 27154 75150 27196
rect 75274 27154 75318 27196
rect 75442 27154 75489 27196
rect 58531 27028 58540 27068
rect 58580 27028 67564 27068
rect 67604 27028 67613 27068
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 16343 26480 16390 26522
rect 16514 26480 16558 26522
rect 16682 26480 16729 26522
rect 16343 26440 16352 26480
rect 16514 26440 16516 26480
rect 16556 26440 16558 26480
rect 16720 26440 16729 26480
rect 16343 26398 16390 26440
rect 16514 26398 16558 26440
rect 16682 26398 16729 26440
rect 28343 26480 28390 26522
rect 28514 26480 28558 26522
rect 28682 26480 28729 26522
rect 28343 26440 28352 26480
rect 28514 26440 28516 26480
rect 28556 26440 28558 26480
rect 28720 26440 28729 26480
rect 28343 26398 28390 26440
rect 28514 26398 28558 26440
rect 28682 26398 28729 26440
rect 40343 26480 40390 26522
rect 40514 26480 40558 26522
rect 40682 26480 40729 26522
rect 40343 26440 40352 26480
rect 40514 26440 40516 26480
rect 40556 26440 40558 26480
rect 40720 26440 40729 26480
rect 40343 26398 40390 26440
rect 40514 26398 40558 26440
rect 40682 26398 40729 26440
rect 52343 26480 52390 26522
rect 52514 26480 52558 26522
rect 52682 26480 52729 26522
rect 64343 26480 64390 26522
rect 64514 26480 64558 26522
rect 64682 26480 64729 26522
rect 52343 26440 52352 26480
rect 52514 26440 52516 26480
rect 52556 26440 52558 26480
rect 52720 26440 52729 26480
rect 52867 26440 52876 26480
rect 52916 26440 54508 26480
rect 54548 26440 54557 26480
rect 64343 26440 64352 26480
rect 64514 26440 64516 26480
rect 64556 26440 64558 26480
rect 64720 26440 64729 26480
rect 52343 26398 52390 26440
rect 52514 26398 52558 26440
rect 52682 26398 52729 26440
rect 64343 26398 64390 26440
rect 64514 26398 64558 26440
rect 64682 26398 64729 26440
rect 76343 26480 76390 26522
rect 76514 26480 76558 26522
rect 76682 26480 76729 26522
rect 76343 26440 76352 26480
rect 76514 26440 76516 26480
rect 76556 26440 76558 26480
rect 76720 26440 76729 26480
rect 76343 26398 76390 26440
rect 76514 26398 76558 26440
rect 76682 26398 76729 26440
rect 56707 26188 56716 26228
rect 56756 26188 60364 26228
rect 60404 26188 60413 26228
rect 43171 26104 43180 26144
rect 43220 26104 56892 26144
rect 56852 26060 56892 26104
rect 40867 26020 40876 26060
rect 40916 26020 56716 26060
rect 56756 26020 56765 26060
rect 56852 26020 60556 26060
rect 60596 26020 60605 26060
rect 38851 25936 38860 25976
rect 38900 25936 58348 25976
rect 58388 25936 58397 25976
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 15103 25724 15150 25766
rect 15274 25724 15318 25766
rect 15442 25724 15489 25766
rect 15103 25684 15112 25724
rect 15274 25684 15276 25724
rect 15316 25684 15318 25724
rect 15480 25684 15489 25724
rect 15103 25642 15150 25684
rect 15274 25642 15318 25684
rect 15442 25642 15489 25684
rect 27103 25724 27150 25766
rect 27274 25724 27318 25766
rect 27442 25724 27489 25766
rect 27103 25684 27112 25724
rect 27274 25684 27276 25724
rect 27316 25684 27318 25724
rect 27480 25684 27489 25724
rect 27103 25642 27150 25684
rect 27274 25642 27318 25684
rect 27442 25642 27489 25684
rect 39103 25724 39150 25766
rect 39274 25724 39318 25766
rect 39442 25724 39489 25766
rect 39103 25684 39112 25724
rect 39274 25684 39276 25724
rect 39316 25684 39318 25724
rect 39480 25684 39489 25724
rect 39103 25642 39150 25684
rect 39274 25642 39318 25684
rect 39442 25642 39489 25684
rect 51103 25724 51150 25766
rect 51274 25724 51318 25766
rect 51442 25724 51489 25766
rect 51103 25684 51112 25724
rect 51274 25684 51276 25724
rect 51316 25684 51318 25724
rect 51480 25684 51489 25724
rect 51103 25642 51150 25684
rect 51274 25642 51318 25684
rect 51442 25642 51489 25684
rect 63103 25724 63150 25766
rect 63274 25724 63318 25766
rect 63442 25724 63489 25766
rect 63103 25684 63112 25724
rect 63274 25684 63276 25724
rect 63316 25684 63318 25724
rect 63480 25684 63489 25724
rect 63103 25642 63150 25684
rect 63274 25642 63318 25684
rect 63442 25642 63489 25684
rect 75103 25724 75150 25766
rect 75274 25724 75318 25766
rect 75442 25724 75489 25766
rect 75103 25684 75112 25724
rect 75274 25684 75276 25724
rect 75316 25684 75318 25724
rect 75480 25684 75489 25724
rect 75103 25642 75150 25684
rect 75274 25642 75318 25684
rect 75442 25642 75489 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 16343 24968 16390 25010
rect 16514 24968 16558 25010
rect 16682 24968 16729 25010
rect 16343 24928 16352 24968
rect 16514 24928 16516 24968
rect 16556 24928 16558 24968
rect 16720 24928 16729 24968
rect 16343 24886 16390 24928
rect 16514 24886 16558 24928
rect 16682 24886 16729 24928
rect 28343 24968 28390 25010
rect 28514 24968 28558 25010
rect 28682 24968 28729 25010
rect 28343 24928 28352 24968
rect 28514 24928 28516 24968
rect 28556 24928 28558 24968
rect 28720 24928 28729 24968
rect 28343 24886 28390 24928
rect 28514 24886 28558 24928
rect 28682 24886 28729 24928
rect 40343 24968 40390 25010
rect 40514 24968 40558 25010
rect 40682 24968 40729 25010
rect 40343 24928 40352 24968
rect 40514 24928 40516 24968
rect 40556 24928 40558 24968
rect 40720 24928 40729 24968
rect 40343 24886 40390 24928
rect 40514 24886 40558 24928
rect 40682 24886 40729 24928
rect 52343 24968 52390 25010
rect 52514 24968 52558 25010
rect 52682 24968 52729 25010
rect 52343 24928 52352 24968
rect 52514 24928 52516 24968
rect 52556 24928 52558 24968
rect 52720 24928 52729 24968
rect 52343 24886 52390 24928
rect 52514 24886 52558 24928
rect 52682 24886 52729 24928
rect 64343 24968 64390 25010
rect 64514 24968 64558 25010
rect 64682 24968 64729 25010
rect 64343 24928 64352 24968
rect 64514 24928 64516 24968
rect 64556 24928 64558 24968
rect 64720 24928 64729 24968
rect 64343 24886 64390 24928
rect 64514 24886 64558 24928
rect 64682 24886 64729 24928
rect 76343 24968 76390 25010
rect 76514 24968 76558 25010
rect 76682 24968 76729 25010
rect 76343 24928 76352 24968
rect 76514 24928 76516 24968
rect 76556 24928 76558 24968
rect 76720 24928 76729 24968
rect 76343 24886 76390 24928
rect 76514 24886 76558 24928
rect 76682 24886 76729 24928
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 15103 24212 15150 24254
rect 15274 24212 15318 24254
rect 15442 24212 15489 24254
rect 15103 24172 15112 24212
rect 15274 24172 15276 24212
rect 15316 24172 15318 24212
rect 15480 24172 15489 24212
rect 15103 24130 15150 24172
rect 15274 24130 15318 24172
rect 15442 24130 15489 24172
rect 27103 24212 27150 24254
rect 27274 24212 27318 24254
rect 27442 24212 27489 24254
rect 27103 24172 27112 24212
rect 27274 24172 27276 24212
rect 27316 24172 27318 24212
rect 27480 24172 27489 24212
rect 27103 24130 27150 24172
rect 27274 24130 27318 24172
rect 27442 24130 27489 24172
rect 39103 24212 39150 24254
rect 39274 24212 39318 24254
rect 39442 24212 39489 24254
rect 39103 24172 39112 24212
rect 39274 24172 39276 24212
rect 39316 24172 39318 24212
rect 39480 24172 39489 24212
rect 39103 24130 39150 24172
rect 39274 24130 39318 24172
rect 39442 24130 39489 24172
rect 51715 23836 51724 23876
rect 51764 23836 54604 23876
rect 54644 23836 54653 23876
rect 78822 23752 79084 23792
rect 79124 23752 79133 23792
rect 48163 23668 48172 23708
rect 48212 23668 55852 23708
rect 55892 23668 55901 23708
rect 48643 23584 48652 23624
rect 48692 23584 54796 23624
rect 54836 23584 54845 23624
rect 50851 23500 50860 23540
rect 50900 23500 56140 23540
rect 56180 23500 56189 23540
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 16343 23456 16390 23498
rect 16514 23456 16558 23498
rect 16682 23456 16729 23498
rect 16343 23416 16352 23456
rect 16514 23416 16516 23456
rect 16556 23416 16558 23456
rect 16720 23416 16729 23456
rect 16343 23374 16390 23416
rect 16514 23374 16558 23416
rect 16682 23374 16729 23416
rect 28343 23456 28390 23498
rect 28514 23456 28558 23498
rect 28682 23456 28729 23498
rect 28343 23416 28352 23456
rect 28514 23416 28516 23456
rect 28556 23416 28558 23456
rect 28720 23416 28729 23456
rect 28343 23374 28390 23416
rect 28514 23374 28558 23416
rect 28682 23374 28729 23416
rect 40343 23456 40390 23498
rect 40514 23456 40558 23498
rect 40682 23456 40729 23498
rect 40343 23416 40352 23456
rect 40514 23416 40516 23456
rect 40556 23416 40558 23456
rect 40720 23416 40729 23456
rect 51619 23416 51628 23456
rect 51668 23416 56812 23456
rect 56852 23416 56861 23456
rect 40343 23374 40390 23416
rect 40514 23374 40558 23416
rect 40682 23374 40729 23416
rect 51811 23332 51820 23372
rect 51860 23332 57292 23372
rect 57332 23332 57676 23372
rect 57716 23332 57725 23372
rect 43180 23248 56812 23288
rect 56852 23248 56861 23288
rect 43180 23204 43220 23248
rect 11683 23164 11692 23204
rect 11732 23164 43220 23204
rect 51523 23164 51532 23204
rect 51572 23164 55660 23204
rect 55700 23164 55709 23204
rect 52579 23080 52588 23120
rect 52628 23080 54412 23120
rect 54452 23080 54461 23120
rect 52483 22828 52492 22868
rect 52532 22828 54700 22868
rect 54740 22828 54749 22868
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 15103 22700 15150 22742
rect 15274 22700 15318 22742
rect 15442 22700 15489 22742
rect 15103 22660 15112 22700
rect 15274 22660 15276 22700
rect 15316 22660 15318 22700
rect 15480 22660 15489 22700
rect 15103 22618 15150 22660
rect 15274 22618 15318 22660
rect 15442 22618 15489 22660
rect 27103 22700 27150 22742
rect 27274 22700 27318 22742
rect 27442 22700 27489 22742
rect 27103 22660 27112 22700
rect 27274 22660 27276 22700
rect 27316 22660 27318 22700
rect 27480 22660 27489 22700
rect 27103 22618 27150 22660
rect 27274 22618 27318 22660
rect 27442 22618 27489 22660
rect 39103 22700 39150 22742
rect 39274 22700 39318 22742
rect 39442 22700 39489 22742
rect 39103 22660 39112 22700
rect 39274 22660 39276 22700
rect 39316 22660 39318 22700
rect 39480 22660 39489 22700
rect 39103 22618 39150 22660
rect 39274 22618 39318 22660
rect 39442 22618 39489 22660
rect 64316 22541 64756 22652
rect 64316 22417 64390 22541
rect 64514 22417 64558 22541
rect 64682 22417 64756 22541
rect 64316 22373 64756 22417
rect 64316 22249 64390 22373
rect 64514 22249 64558 22373
rect 64682 22249 64756 22373
rect 64316 22205 64756 22249
rect 64316 22081 64390 22205
rect 64514 22081 64558 22205
rect 64682 22081 64756 22205
rect 64316 22037 64756 22081
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 16343 21944 16390 21986
rect 16514 21944 16558 21986
rect 16682 21944 16729 21986
rect 16343 21904 16352 21944
rect 16514 21904 16516 21944
rect 16556 21904 16558 21944
rect 16720 21904 16729 21944
rect 16343 21862 16390 21904
rect 16514 21862 16558 21904
rect 16682 21862 16729 21904
rect 28343 21944 28390 21986
rect 28514 21944 28558 21986
rect 28682 21944 28729 21986
rect 28343 21904 28352 21944
rect 28514 21904 28516 21944
rect 28556 21904 28558 21944
rect 28720 21904 28729 21944
rect 28343 21862 28390 21904
rect 28514 21862 28558 21904
rect 28682 21862 28729 21904
rect 40343 21944 40390 21986
rect 40514 21944 40558 21986
rect 40682 21944 40729 21986
rect 40343 21904 40352 21944
rect 40514 21904 40516 21944
rect 40556 21904 40558 21944
rect 40720 21904 40729 21944
rect 40343 21862 40390 21904
rect 40514 21862 40558 21904
rect 40682 21862 40729 21904
rect 64316 21913 64390 22037
rect 64514 21913 64558 22037
rect 64682 21913 64756 22037
rect 64316 21869 64756 21913
rect 64316 21745 64390 21869
rect 64514 21745 64558 21869
rect 64682 21745 64756 21869
rect 64316 21701 64756 21745
rect 64316 21577 64390 21701
rect 64514 21577 64558 21701
rect 64682 21577 64756 21701
rect 64316 21533 64756 21577
rect 64316 21409 64390 21533
rect 64514 21409 64558 21533
rect 64682 21409 64756 21533
rect 64316 21365 64756 21409
rect 64316 21241 64390 21365
rect 64514 21241 64558 21365
rect 64682 21241 64756 21365
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 15103 21188 15150 21230
rect 15274 21188 15318 21230
rect 15442 21188 15489 21230
rect 15103 21148 15112 21188
rect 15274 21148 15276 21188
rect 15316 21148 15318 21188
rect 15480 21148 15489 21188
rect 15103 21106 15150 21148
rect 15274 21106 15318 21148
rect 15442 21106 15489 21148
rect 27103 21188 27150 21230
rect 27274 21188 27318 21230
rect 27442 21188 27489 21230
rect 27103 21148 27112 21188
rect 27274 21148 27276 21188
rect 27316 21148 27318 21188
rect 27480 21148 27489 21188
rect 27103 21106 27150 21148
rect 27274 21106 27318 21148
rect 27442 21106 27489 21148
rect 39103 21188 39150 21230
rect 39274 21188 39318 21230
rect 39442 21188 39489 21230
rect 39103 21148 39112 21188
rect 39274 21148 39276 21188
rect 39316 21148 39318 21188
rect 39480 21148 39489 21188
rect 39103 21106 39150 21148
rect 39274 21106 39318 21148
rect 39442 21106 39489 21148
rect 64316 21197 64756 21241
rect 64316 21073 64390 21197
rect 64514 21073 64558 21197
rect 64682 21073 64756 21197
rect 64316 21029 64756 21073
rect 64316 20905 64390 21029
rect 64514 20905 64558 21029
rect 64682 20905 64756 21029
rect 64316 20861 64756 20905
rect 64316 20737 64390 20861
rect 64514 20737 64558 20861
rect 64682 20737 64756 20861
rect 64316 20693 64756 20737
rect 64316 20569 64390 20693
rect 64514 20569 64558 20693
rect 64682 20569 64756 20693
rect 64316 20525 64756 20569
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 16343 20432 16390 20474
rect 16514 20432 16558 20474
rect 16682 20432 16729 20474
rect 16343 20392 16352 20432
rect 16514 20392 16516 20432
rect 16556 20392 16558 20432
rect 16720 20392 16729 20432
rect 16343 20350 16390 20392
rect 16514 20350 16558 20392
rect 16682 20350 16729 20392
rect 28343 20432 28390 20474
rect 28514 20432 28558 20474
rect 28682 20432 28729 20474
rect 28343 20392 28352 20432
rect 28514 20392 28516 20432
rect 28556 20392 28558 20432
rect 28720 20392 28729 20432
rect 28343 20350 28390 20392
rect 28514 20350 28558 20392
rect 28682 20350 28729 20392
rect 40343 20432 40390 20474
rect 40514 20432 40558 20474
rect 40682 20432 40729 20474
rect 40343 20392 40352 20432
rect 40514 20392 40516 20432
rect 40556 20392 40558 20432
rect 40720 20392 40729 20432
rect 40343 20350 40390 20392
rect 40514 20350 40558 20392
rect 40682 20350 40729 20392
rect 64316 20401 64390 20525
rect 64514 20401 64558 20525
rect 64682 20401 64756 20525
rect 64316 20290 64756 20401
rect 76316 22541 76756 22652
rect 76316 22417 76390 22541
rect 76514 22417 76558 22541
rect 76682 22417 76756 22541
rect 76316 22373 76756 22417
rect 76316 22249 76390 22373
rect 76514 22249 76558 22373
rect 76682 22249 76756 22373
rect 76316 22205 76756 22249
rect 76316 22081 76390 22205
rect 76514 22081 76558 22205
rect 76682 22081 76756 22205
rect 76316 22037 76756 22081
rect 76316 21913 76390 22037
rect 76514 21913 76558 22037
rect 76682 21913 76756 22037
rect 76316 21869 76756 21913
rect 76316 21745 76390 21869
rect 76514 21745 76558 21869
rect 76682 21745 76756 21869
rect 76316 21701 76756 21745
rect 76316 21577 76390 21701
rect 76514 21577 76558 21701
rect 76682 21577 76756 21701
rect 76316 21533 76756 21577
rect 76316 21409 76390 21533
rect 76514 21409 76558 21533
rect 76682 21409 76756 21533
rect 76316 21365 76756 21409
rect 76316 21241 76390 21365
rect 76514 21241 76558 21365
rect 76682 21241 76756 21365
rect 76316 21197 76756 21241
rect 76316 21073 76390 21197
rect 76514 21073 76558 21197
rect 76682 21073 76756 21197
rect 76316 21029 76756 21073
rect 76316 20905 76390 21029
rect 76514 20905 76558 21029
rect 76682 20905 76756 21029
rect 76316 20861 76756 20905
rect 76316 20737 76390 20861
rect 76514 20737 76558 20861
rect 76682 20737 76756 20861
rect 76316 20693 76756 20737
rect 76316 20569 76390 20693
rect 76514 20569 76558 20693
rect 76682 20569 76756 20693
rect 76316 20525 76756 20569
rect 76316 20401 76390 20525
rect 76514 20401 76558 20525
rect 76682 20401 76756 20525
rect 76316 20290 76756 20401
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 15103 19676 15150 19718
rect 15274 19676 15318 19718
rect 15442 19676 15489 19718
rect 15103 19636 15112 19676
rect 15274 19636 15276 19676
rect 15316 19636 15318 19676
rect 15480 19636 15489 19676
rect 15103 19594 15150 19636
rect 15274 19594 15318 19636
rect 15442 19594 15489 19636
rect 27103 19676 27150 19718
rect 27274 19676 27318 19718
rect 27442 19676 27489 19718
rect 27103 19636 27112 19676
rect 27274 19636 27276 19676
rect 27316 19636 27318 19676
rect 27480 19636 27489 19676
rect 27103 19594 27150 19636
rect 27274 19594 27318 19636
rect 27442 19594 27489 19636
rect 39103 19676 39150 19718
rect 39274 19676 39318 19718
rect 39442 19676 39489 19718
rect 39103 19636 39112 19676
rect 39274 19636 39276 19676
rect 39316 19636 39318 19676
rect 39480 19636 39489 19676
rect 39103 19594 39150 19636
rect 39274 19594 39318 19636
rect 39442 19594 39489 19636
rect 63076 19665 63516 19776
rect 63076 19541 63150 19665
rect 63274 19541 63318 19665
rect 63442 19541 63516 19665
rect 63076 19497 63516 19541
rect 63076 19373 63150 19497
rect 63274 19373 63318 19497
rect 63442 19373 63516 19497
rect 63076 19329 63516 19373
rect 63076 19205 63150 19329
rect 63274 19205 63318 19329
rect 63442 19205 63516 19329
rect 63076 19161 63516 19205
rect 63076 19037 63150 19161
rect 63274 19037 63318 19161
rect 63442 19037 63516 19161
rect 63076 18993 63516 19037
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 16343 18920 16390 18962
rect 16514 18920 16558 18962
rect 16682 18920 16729 18962
rect 16343 18880 16352 18920
rect 16514 18880 16516 18920
rect 16556 18880 16558 18920
rect 16720 18880 16729 18920
rect 16343 18838 16390 18880
rect 16514 18838 16558 18880
rect 16682 18838 16729 18880
rect 28343 18920 28390 18962
rect 28514 18920 28558 18962
rect 28682 18920 28729 18962
rect 28343 18880 28352 18920
rect 28514 18880 28516 18920
rect 28556 18880 28558 18920
rect 28720 18880 28729 18920
rect 28343 18838 28390 18880
rect 28514 18838 28558 18880
rect 28682 18838 28729 18880
rect 40343 18920 40390 18962
rect 40514 18920 40558 18962
rect 40682 18920 40729 18962
rect 40343 18880 40352 18920
rect 40514 18880 40516 18920
rect 40556 18880 40558 18920
rect 40720 18880 40729 18920
rect 40343 18838 40390 18880
rect 40514 18838 40558 18880
rect 40682 18838 40729 18880
rect 63076 18869 63150 18993
rect 63274 18869 63318 18993
rect 63442 18869 63516 18993
rect 63076 18825 63516 18869
rect 63076 18701 63150 18825
rect 63274 18701 63318 18825
rect 63442 18701 63516 18825
rect 63076 18657 63516 18701
rect 63076 18533 63150 18657
rect 63274 18533 63318 18657
rect 63442 18533 63516 18657
rect 43075 18460 43084 18500
rect 43124 18460 51340 18500
rect 51380 18460 51389 18500
rect 63076 18489 63516 18533
rect 63076 18365 63150 18489
rect 63274 18365 63318 18489
rect 63442 18365 63516 18489
rect 35395 18292 35404 18332
rect 35444 18292 50380 18332
rect 50420 18292 50429 18332
rect 63076 18321 63516 18365
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 15103 18164 15150 18206
rect 15274 18164 15318 18206
rect 15442 18164 15489 18206
rect 15103 18124 15112 18164
rect 15274 18124 15276 18164
rect 15316 18124 15318 18164
rect 15480 18124 15489 18164
rect 15103 18082 15150 18124
rect 15274 18082 15318 18124
rect 15442 18082 15489 18124
rect 27103 18164 27150 18206
rect 27274 18164 27318 18206
rect 27442 18164 27489 18206
rect 27103 18124 27112 18164
rect 27274 18124 27276 18164
rect 27316 18124 27318 18164
rect 27480 18124 27489 18164
rect 27103 18082 27150 18124
rect 27274 18082 27318 18124
rect 27442 18082 27489 18124
rect 39103 18164 39150 18206
rect 39274 18164 39318 18206
rect 39442 18164 39489 18206
rect 39103 18124 39112 18164
rect 39274 18124 39276 18164
rect 39316 18124 39318 18164
rect 39480 18124 39489 18164
rect 39103 18082 39150 18124
rect 39274 18082 39318 18124
rect 39442 18082 39489 18124
rect 63076 18197 63150 18321
rect 63274 18197 63318 18321
rect 63442 18197 63516 18321
rect 63076 18153 63516 18197
rect 63076 18029 63150 18153
rect 63274 18029 63318 18153
rect 63442 18029 63516 18153
rect 63076 17985 63516 18029
rect 63076 17861 63150 17985
rect 63274 17861 63318 17985
rect 63442 17861 63516 17985
rect 63076 17817 63516 17861
rect 63076 17693 63150 17817
rect 63274 17693 63318 17817
rect 63442 17693 63516 17817
rect 63076 17649 63516 17693
rect 25507 17536 25516 17576
rect 25556 17536 52300 17576
rect 52340 17536 52349 17576
rect 63076 17525 63150 17649
rect 63274 17525 63318 17649
rect 63442 17525 63516 17649
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 16343 17408 16390 17450
rect 16514 17408 16558 17450
rect 16682 17408 16729 17450
rect 16343 17368 16352 17408
rect 16514 17368 16516 17408
rect 16556 17368 16558 17408
rect 16720 17368 16729 17408
rect 16343 17326 16390 17368
rect 16514 17326 16558 17368
rect 16682 17326 16729 17368
rect 28343 17408 28390 17450
rect 28514 17408 28558 17450
rect 28682 17408 28729 17450
rect 28343 17368 28352 17408
rect 28514 17368 28516 17408
rect 28556 17368 28558 17408
rect 28720 17368 28729 17408
rect 28343 17326 28390 17368
rect 28514 17326 28558 17368
rect 28682 17326 28729 17368
rect 40343 17408 40390 17450
rect 40514 17408 40558 17450
rect 40682 17408 40729 17450
rect 63076 17414 63516 17525
rect 75076 19665 75516 19776
rect 75076 19541 75150 19665
rect 75274 19541 75318 19665
rect 75442 19541 75516 19665
rect 75076 19497 75516 19541
rect 75076 19373 75150 19497
rect 75274 19373 75318 19497
rect 75442 19373 75516 19497
rect 75076 19329 75516 19373
rect 75076 19205 75150 19329
rect 75274 19205 75318 19329
rect 75442 19205 75516 19329
rect 75076 19161 75516 19205
rect 75076 19037 75150 19161
rect 75274 19037 75318 19161
rect 75442 19037 75516 19161
rect 75076 18993 75516 19037
rect 75076 18869 75150 18993
rect 75274 18869 75318 18993
rect 75442 18869 75516 18993
rect 75076 18825 75516 18869
rect 75076 18701 75150 18825
rect 75274 18701 75318 18825
rect 75442 18701 75516 18825
rect 75076 18657 75516 18701
rect 75076 18533 75150 18657
rect 75274 18533 75318 18657
rect 75442 18533 75516 18657
rect 75076 18489 75516 18533
rect 75076 18365 75150 18489
rect 75274 18365 75318 18489
rect 75442 18365 75516 18489
rect 75076 18321 75516 18365
rect 75076 18197 75150 18321
rect 75274 18197 75318 18321
rect 75442 18197 75516 18321
rect 75076 18153 75516 18197
rect 75076 18029 75150 18153
rect 75274 18029 75318 18153
rect 75442 18029 75516 18153
rect 75076 17985 75516 18029
rect 75076 17861 75150 17985
rect 75274 17861 75318 17985
rect 75442 17861 75516 17985
rect 75076 17817 75516 17861
rect 75076 17693 75150 17817
rect 75274 17693 75318 17817
rect 75442 17693 75516 17817
rect 75076 17649 75516 17693
rect 75076 17525 75150 17649
rect 75274 17525 75318 17649
rect 75442 17525 75516 17649
rect 75076 17414 75516 17525
rect 40343 17368 40352 17408
rect 40514 17368 40516 17408
rect 40556 17368 40558 17408
rect 40720 17368 40729 17408
rect 40343 17326 40390 17368
rect 40514 17326 40558 17368
rect 40682 17326 40729 17368
rect 50371 17200 50380 17240
rect 50420 17200 55084 17240
rect 55124 17200 55133 17240
rect 52291 17116 52300 17156
rect 52340 17116 52780 17156
rect 52820 17116 52829 17156
rect 52579 17032 52588 17072
rect 52628 17032 78892 17072
rect 78932 17032 78941 17072
rect 32803 16948 32812 16988
rect 32852 16948 54700 16988
rect 54740 16948 54749 16988
rect 36643 16864 36652 16904
rect 36692 16864 58252 16904
rect 58292 16864 58301 16904
rect 29635 16780 29644 16820
rect 29684 16780 51916 16820
rect 51956 16780 54316 16820
rect 54356 16780 54365 16820
rect 39715 16696 39724 16736
rect 39764 16696 57868 16736
rect 57908 16696 57917 16736
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 15103 16652 15150 16694
rect 15274 16652 15318 16694
rect 15442 16652 15489 16694
rect 15103 16612 15112 16652
rect 15274 16612 15276 16652
rect 15316 16612 15318 16652
rect 15480 16612 15489 16652
rect 15103 16570 15150 16612
rect 15274 16570 15318 16612
rect 15442 16570 15489 16612
rect 27103 16652 27150 16694
rect 27274 16652 27318 16694
rect 27442 16652 27489 16694
rect 27103 16612 27112 16652
rect 27274 16612 27276 16652
rect 27316 16612 27318 16652
rect 27480 16612 27489 16652
rect 27103 16570 27150 16612
rect 27274 16570 27318 16612
rect 27442 16570 27489 16612
rect 39103 16652 39150 16694
rect 39274 16652 39318 16694
rect 39442 16652 39489 16694
rect 39103 16612 39112 16652
rect 39274 16612 39276 16652
rect 39316 16612 39318 16652
rect 39480 16612 39489 16652
rect 39103 16570 39150 16612
rect 39274 16570 39318 16612
rect 39442 16570 39489 16612
rect 52003 16276 52012 16316
rect 52052 16276 61708 16316
rect 61748 16276 61757 16316
rect 51811 16192 51820 16232
rect 51860 16192 64972 16232
rect 65012 16192 65021 16232
rect 78822 16192 78892 16232
rect 78932 16192 78941 16232
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 16343 15896 16390 15938
rect 16514 15896 16558 15938
rect 16682 15896 16729 15938
rect 16343 15856 16352 15896
rect 16514 15856 16516 15896
rect 16556 15856 16558 15896
rect 16720 15856 16729 15896
rect 16343 15814 16390 15856
rect 16514 15814 16558 15856
rect 16682 15814 16729 15856
rect 28343 15896 28390 15938
rect 28514 15896 28558 15938
rect 28682 15896 28729 15938
rect 28343 15856 28352 15896
rect 28514 15856 28516 15896
rect 28556 15856 28558 15896
rect 28720 15856 28729 15896
rect 28343 15814 28390 15856
rect 28514 15814 28558 15856
rect 28682 15814 28729 15856
rect 40343 15896 40390 15938
rect 40514 15896 40558 15938
rect 40682 15896 40729 15938
rect 40343 15856 40352 15896
rect 40514 15856 40516 15896
rect 40556 15856 40558 15896
rect 40720 15856 40729 15896
rect 40343 15814 40390 15856
rect 40514 15814 40558 15856
rect 40682 15814 40729 15856
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 15103 15140 15150 15182
rect 15274 15140 15318 15182
rect 15442 15140 15489 15182
rect 15103 15100 15112 15140
rect 15274 15100 15276 15140
rect 15316 15100 15318 15140
rect 15480 15100 15489 15140
rect 15103 15058 15150 15100
rect 15274 15058 15318 15100
rect 15442 15058 15489 15100
rect 27103 15140 27150 15182
rect 27274 15140 27318 15182
rect 27442 15140 27489 15182
rect 27103 15100 27112 15140
rect 27274 15100 27276 15140
rect 27316 15100 27318 15140
rect 27480 15100 27489 15140
rect 27103 15058 27150 15100
rect 27274 15058 27318 15100
rect 27442 15058 27489 15100
rect 39103 15140 39150 15182
rect 39274 15140 39318 15182
rect 39442 15140 39489 15182
rect 39103 15100 39112 15140
rect 39274 15100 39276 15140
rect 39316 15100 39318 15140
rect 39480 15100 39489 15140
rect 39103 15058 39150 15100
rect 39274 15058 39318 15100
rect 39442 15058 39489 15100
rect 51103 15140 51150 15182
rect 51274 15140 51318 15182
rect 51442 15140 51489 15182
rect 51103 15100 51112 15140
rect 51274 15100 51276 15140
rect 51316 15100 51318 15140
rect 51480 15100 51489 15140
rect 51103 15058 51150 15100
rect 51274 15058 51318 15100
rect 51442 15058 51489 15100
rect 63103 15140 63150 15182
rect 63274 15140 63318 15182
rect 63442 15140 63489 15182
rect 63103 15100 63112 15140
rect 63274 15100 63276 15140
rect 63316 15100 63318 15140
rect 63480 15100 63489 15140
rect 63103 15058 63150 15100
rect 63274 15058 63318 15100
rect 63442 15058 63489 15100
rect 75103 15140 75150 15182
rect 75274 15140 75318 15182
rect 75442 15140 75489 15182
rect 75103 15100 75112 15140
rect 75274 15100 75276 15140
rect 75316 15100 75318 15140
rect 75480 15100 75489 15140
rect 75103 15058 75150 15100
rect 75274 15058 75318 15100
rect 75442 15058 75489 15100
rect 52867 14932 52876 14972
rect 52916 14932 61900 14972
rect 61940 14932 61949 14972
rect 53059 14848 53068 14888
rect 53108 14848 60748 14888
rect 60788 14848 60797 14888
rect 52099 14764 52108 14804
rect 52148 14764 58924 14804
rect 58964 14764 67180 14804
rect 67220 14764 67229 14804
rect 32323 14512 32332 14552
rect 32372 14512 58540 14552
rect 58580 14512 58589 14552
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 16343 14384 16390 14426
rect 16514 14384 16558 14426
rect 16682 14384 16729 14426
rect 16343 14344 16352 14384
rect 16514 14344 16516 14384
rect 16556 14344 16558 14384
rect 16720 14344 16729 14384
rect 16343 14302 16390 14344
rect 16514 14302 16558 14344
rect 16682 14302 16729 14344
rect 28343 14384 28390 14426
rect 28514 14384 28558 14426
rect 28682 14384 28729 14426
rect 28343 14344 28352 14384
rect 28514 14344 28516 14384
rect 28556 14344 28558 14384
rect 28720 14344 28729 14384
rect 28343 14302 28390 14344
rect 28514 14302 28558 14344
rect 28682 14302 28729 14344
rect 40343 14384 40390 14426
rect 40514 14384 40558 14426
rect 40682 14384 40729 14426
rect 40343 14344 40352 14384
rect 40514 14344 40516 14384
rect 40556 14344 40558 14384
rect 40720 14344 40729 14384
rect 40343 14302 40390 14344
rect 40514 14302 40558 14344
rect 40682 14302 40729 14344
rect 52343 14384 52390 14426
rect 52514 14384 52558 14426
rect 52682 14384 52729 14426
rect 52343 14344 52352 14384
rect 52514 14344 52516 14384
rect 52556 14344 52558 14384
rect 52720 14344 52729 14384
rect 52343 14302 52390 14344
rect 52514 14302 52558 14344
rect 52682 14302 52729 14344
rect 64343 14384 64390 14426
rect 64514 14384 64558 14426
rect 64682 14384 64729 14426
rect 64343 14344 64352 14384
rect 64514 14344 64516 14384
rect 64556 14344 64558 14384
rect 64720 14344 64729 14384
rect 64343 14302 64390 14344
rect 64514 14302 64558 14344
rect 64682 14302 64729 14344
rect 76343 14384 76390 14426
rect 76514 14384 76558 14426
rect 76682 14384 76729 14426
rect 76343 14344 76352 14384
rect 76514 14344 76516 14384
rect 76556 14344 76558 14384
rect 76720 14344 76729 14384
rect 76343 14302 76390 14344
rect 76514 14302 76558 14344
rect 76682 14302 76729 14344
rect 57859 13924 57868 13964
rect 57908 13924 69196 13964
rect 69236 13924 69245 13964
rect 51907 13840 51916 13880
rect 51956 13840 57772 13880
rect 57812 13840 57821 13880
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 15103 13628 15150 13670
rect 15274 13628 15318 13670
rect 15442 13628 15489 13670
rect 15103 13588 15112 13628
rect 15274 13588 15276 13628
rect 15316 13588 15318 13628
rect 15480 13588 15489 13628
rect 15103 13546 15150 13588
rect 15274 13546 15318 13588
rect 15442 13546 15489 13588
rect 27103 13628 27150 13670
rect 27274 13628 27318 13670
rect 27442 13628 27489 13670
rect 27103 13588 27112 13628
rect 27274 13588 27276 13628
rect 27316 13588 27318 13628
rect 27480 13588 27489 13628
rect 27103 13546 27150 13588
rect 27274 13546 27318 13588
rect 27442 13546 27489 13588
rect 39103 13628 39150 13670
rect 39274 13628 39318 13670
rect 39442 13628 39489 13670
rect 39103 13588 39112 13628
rect 39274 13588 39276 13628
rect 39316 13588 39318 13628
rect 39480 13588 39489 13628
rect 39103 13546 39150 13588
rect 39274 13546 39318 13588
rect 39442 13546 39489 13588
rect 51103 13628 51150 13670
rect 51274 13628 51318 13670
rect 51442 13628 51489 13670
rect 51103 13588 51112 13628
rect 51274 13588 51276 13628
rect 51316 13588 51318 13628
rect 51480 13588 51489 13628
rect 51103 13546 51150 13588
rect 51274 13546 51318 13588
rect 51442 13546 51489 13588
rect 63103 13628 63150 13670
rect 63274 13628 63318 13670
rect 63442 13628 63489 13670
rect 63103 13588 63112 13628
rect 63274 13588 63276 13628
rect 63316 13588 63318 13628
rect 63480 13588 63489 13628
rect 63103 13546 63150 13588
rect 63274 13546 63318 13588
rect 63442 13546 63489 13588
rect 75103 13628 75150 13670
rect 75274 13628 75318 13670
rect 75442 13628 75489 13670
rect 75103 13588 75112 13628
rect 75274 13588 75276 13628
rect 75316 13588 75318 13628
rect 75480 13588 75489 13628
rect 75103 13546 75150 13588
rect 75274 13546 75318 13588
rect 75442 13546 75489 13588
rect 52963 13000 52972 13040
rect 53012 13000 57868 13040
rect 57908 13000 57917 13040
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 16343 12872 16390 12914
rect 16514 12872 16558 12914
rect 16682 12872 16729 12914
rect 16343 12832 16352 12872
rect 16514 12832 16516 12872
rect 16556 12832 16558 12872
rect 16720 12832 16729 12872
rect 16343 12790 16390 12832
rect 16514 12790 16558 12832
rect 16682 12790 16729 12832
rect 28343 12872 28390 12914
rect 28514 12872 28558 12914
rect 28682 12872 28729 12914
rect 28343 12832 28352 12872
rect 28514 12832 28516 12872
rect 28556 12832 28558 12872
rect 28720 12832 28729 12872
rect 28343 12790 28390 12832
rect 28514 12790 28558 12832
rect 28682 12790 28729 12832
rect 40343 12872 40390 12914
rect 40514 12872 40558 12914
rect 40682 12872 40729 12914
rect 40343 12832 40352 12872
rect 40514 12832 40516 12872
rect 40556 12832 40558 12872
rect 40720 12832 40729 12872
rect 40343 12790 40390 12832
rect 40514 12790 40558 12832
rect 40682 12790 40729 12832
rect 52343 12872 52390 12914
rect 52514 12872 52558 12914
rect 52682 12872 52729 12914
rect 52343 12832 52352 12872
rect 52514 12832 52516 12872
rect 52556 12832 52558 12872
rect 52720 12832 52729 12872
rect 52343 12790 52390 12832
rect 52514 12790 52558 12832
rect 52682 12790 52729 12832
rect 64343 12872 64390 12914
rect 64514 12872 64558 12914
rect 64682 12872 64729 12914
rect 64343 12832 64352 12872
rect 64514 12832 64516 12872
rect 64556 12832 64558 12872
rect 64720 12832 64729 12872
rect 64343 12790 64390 12832
rect 64514 12790 64558 12832
rect 64682 12790 64729 12832
rect 76343 12872 76390 12914
rect 76514 12872 76558 12914
rect 76682 12872 76729 12914
rect 76343 12832 76352 12872
rect 76514 12832 76516 12872
rect 76556 12832 76558 12872
rect 76720 12832 76729 12872
rect 76343 12790 76390 12832
rect 76514 12790 76558 12832
rect 76682 12790 76729 12832
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 15103 12116 15150 12158
rect 15274 12116 15318 12158
rect 15442 12116 15489 12158
rect 15103 12076 15112 12116
rect 15274 12076 15276 12116
rect 15316 12076 15318 12116
rect 15480 12076 15489 12116
rect 15103 12034 15150 12076
rect 15274 12034 15318 12076
rect 15442 12034 15489 12076
rect 27103 12116 27150 12158
rect 27274 12116 27318 12158
rect 27442 12116 27489 12158
rect 27103 12076 27112 12116
rect 27274 12076 27276 12116
rect 27316 12076 27318 12116
rect 27480 12076 27489 12116
rect 27103 12034 27150 12076
rect 27274 12034 27318 12076
rect 27442 12034 27489 12076
rect 39103 12116 39150 12158
rect 39274 12116 39318 12158
rect 39442 12116 39489 12158
rect 39103 12076 39112 12116
rect 39274 12076 39276 12116
rect 39316 12076 39318 12116
rect 39480 12076 39489 12116
rect 39103 12034 39150 12076
rect 39274 12034 39318 12076
rect 39442 12034 39489 12076
rect 51103 12116 51150 12158
rect 51274 12116 51318 12158
rect 51442 12116 51489 12158
rect 51103 12076 51112 12116
rect 51274 12076 51276 12116
rect 51316 12076 51318 12116
rect 51480 12076 51489 12116
rect 51103 12034 51150 12076
rect 51274 12034 51318 12076
rect 51442 12034 51489 12076
rect 63103 12116 63150 12158
rect 63274 12116 63318 12158
rect 63442 12116 63489 12158
rect 63103 12076 63112 12116
rect 63274 12076 63276 12116
rect 63316 12076 63318 12116
rect 63480 12076 63489 12116
rect 63103 12034 63150 12076
rect 63274 12034 63318 12076
rect 63442 12034 63489 12076
rect 75103 12116 75150 12158
rect 75274 12116 75318 12158
rect 75442 12116 75489 12158
rect 75103 12076 75112 12116
rect 75274 12076 75276 12116
rect 75316 12076 75318 12116
rect 75480 12076 75489 12116
rect 75103 12034 75150 12076
rect 75274 12034 75318 12076
rect 75442 12034 75489 12076
rect 70531 11572 70540 11612
rect 70580 11572 76204 11612
rect 76244 11572 76396 11612
rect 76436 11572 76445 11612
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 16343 11360 16390 11402
rect 16514 11360 16558 11402
rect 16682 11360 16729 11402
rect 16343 11320 16352 11360
rect 16514 11320 16516 11360
rect 16556 11320 16558 11360
rect 16720 11320 16729 11360
rect 16343 11278 16390 11320
rect 16514 11278 16558 11320
rect 16682 11278 16729 11320
rect 28343 11360 28390 11402
rect 28514 11360 28558 11402
rect 28682 11360 28729 11402
rect 28343 11320 28352 11360
rect 28514 11320 28516 11360
rect 28556 11320 28558 11360
rect 28720 11320 28729 11360
rect 28343 11278 28390 11320
rect 28514 11278 28558 11320
rect 28682 11278 28729 11320
rect 40343 11360 40390 11402
rect 40514 11360 40558 11402
rect 40682 11360 40729 11402
rect 40343 11320 40352 11360
rect 40514 11320 40516 11360
rect 40556 11320 40558 11360
rect 40720 11320 40729 11360
rect 40343 11278 40390 11320
rect 40514 11278 40558 11320
rect 40682 11278 40729 11320
rect 52343 11360 52390 11402
rect 52514 11360 52558 11402
rect 52682 11360 52729 11402
rect 52343 11320 52352 11360
rect 52514 11320 52516 11360
rect 52556 11320 52558 11360
rect 52720 11320 52729 11360
rect 52343 11278 52390 11320
rect 52514 11278 52558 11320
rect 52682 11278 52729 11320
rect 64343 11360 64390 11402
rect 64514 11360 64558 11402
rect 64682 11360 64729 11402
rect 64343 11320 64352 11360
rect 64514 11320 64516 11360
rect 64556 11320 64558 11360
rect 64720 11320 64729 11360
rect 64343 11278 64390 11320
rect 64514 11278 64558 11320
rect 64682 11278 64729 11320
rect 76343 11360 76390 11402
rect 76514 11360 76558 11402
rect 76682 11360 76729 11402
rect 76343 11320 76352 11360
rect 76514 11320 76516 11360
rect 76556 11320 76558 11360
rect 76720 11320 76729 11360
rect 76343 11278 76390 11320
rect 76514 11278 76558 11320
rect 76682 11278 76729 11320
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 15103 10604 15150 10646
rect 15274 10604 15318 10646
rect 15442 10604 15489 10646
rect 15103 10564 15112 10604
rect 15274 10564 15276 10604
rect 15316 10564 15318 10604
rect 15480 10564 15489 10604
rect 15103 10522 15150 10564
rect 15274 10522 15318 10564
rect 15442 10522 15489 10564
rect 27103 10604 27150 10646
rect 27274 10604 27318 10646
rect 27442 10604 27489 10646
rect 27103 10564 27112 10604
rect 27274 10564 27276 10604
rect 27316 10564 27318 10604
rect 27480 10564 27489 10604
rect 27103 10522 27150 10564
rect 27274 10522 27318 10564
rect 27442 10522 27489 10564
rect 39103 10604 39150 10646
rect 39274 10604 39318 10646
rect 39442 10604 39489 10646
rect 39103 10564 39112 10604
rect 39274 10564 39276 10604
rect 39316 10564 39318 10604
rect 39480 10564 39489 10604
rect 39103 10522 39150 10564
rect 39274 10522 39318 10564
rect 39442 10522 39489 10564
rect 51103 10604 51150 10646
rect 51274 10604 51318 10646
rect 51442 10604 51489 10646
rect 51103 10564 51112 10604
rect 51274 10564 51276 10604
rect 51316 10564 51318 10604
rect 51480 10564 51489 10604
rect 51103 10522 51150 10564
rect 51274 10522 51318 10564
rect 51442 10522 51489 10564
rect 63103 10604 63150 10646
rect 63274 10604 63318 10646
rect 63442 10604 63489 10646
rect 63103 10564 63112 10604
rect 63274 10564 63276 10604
rect 63316 10564 63318 10604
rect 63480 10564 63489 10604
rect 63103 10522 63150 10564
rect 63274 10522 63318 10564
rect 63442 10522 63489 10564
rect 75103 10604 75150 10646
rect 75274 10604 75318 10646
rect 75442 10604 75489 10646
rect 75103 10564 75112 10604
rect 75274 10564 75276 10604
rect 75316 10564 75318 10604
rect 75480 10564 75489 10604
rect 75103 10522 75150 10564
rect 75274 10522 75318 10564
rect 75442 10522 75489 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 16343 9848 16390 9890
rect 16514 9848 16558 9890
rect 16682 9848 16729 9890
rect 16343 9808 16352 9848
rect 16514 9808 16516 9848
rect 16556 9808 16558 9848
rect 16720 9808 16729 9848
rect 16343 9766 16390 9808
rect 16514 9766 16558 9808
rect 16682 9766 16729 9808
rect 28343 9848 28390 9890
rect 28514 9848 28558 9890
rect 28682 9848 28729 9890
rect 28343 9808 28352 9848
rect 28514 9808 28516 9848
rect 28556 9808 28558 9848
rect 28720 9808 28729 9848
rect 28343 9766 28390 9808
rect 28514 9766 28558 9808
rect 28682 9766 28729 9808
rect 40343 9848 40390 9890
rect 40514 9848 40558 9890
rect 40682 9848 40729 9890
rect 40343 9808 40352 9848
rect 40514 9808 40516 9848
rect 40556 9808 40558 9848
rect 40720 9808 40729 9848
rect 40343 9766 40390 9808
rect 40514 9766 40558 9808
rect 40682 9766 40729 9808
rect 52343 9848 52390 9890
rect 52514 9848 52558 9890
rect 52682 9848 52729 9890
rect 52343 9808 52352 9848
rect 52514 9808 52516 9848
rect 52556 9808 52558 9848
rect 52720 9808 52729 9848
rect 52343 9766 52390 9808
rect 52514 9766 52558 9808
rect 52682 9766 52729 9808
rect 64343 9848 64390 9890
rect 64514 9848 64558 9890
rect 64682 9848 64729 9890
rect 64343 9808 64352 9848
rect 64514 9808 64516 9848
rect 64556 9808 64558 9848
rect 64720 9808 64729 9848
rect 64343 9766 64390 9808
rect 64514 9766 64558 9808
rect 64682 9766 64729 9808
rect 76343 9848 76390 9890
rect 76514 9848 76558 9890
rect 76682 9848 76729 9890
rect 76343 9808 76352 9848
rect 76514 9808 76516 9848
rect 76556 9808 76558 9848
rect 76720 9808 76729 9848
rect 76343 9766 76390 9808
rect 76514 9766 76558 9808
rect 76682 9766 76729 9808
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 15103 9092 15150 9134
rect 15274 9092 15318 9134
rect 15442 9092 15489 9134
rect 15103 9052 15112 9092
rect 15274 9052 15276 9092
rect 15316 9052 15318 9092
rect 15480 9052 15489 9092
rect 15103 9010 15150 9052
rect 15274 9010 15318 9052
rect 15442 9010 15489 9052
rect 27103 9092 27150 9134
rect 27274 9092 27318 9134
rect 27442 9092 27489 9134
rect 27103 9052 27112 9092
rect 27274 9052 27276 9092
rect 27316 9052 27318 9092
rect 27480 9052 27489 9092
rect 27103 9010 27150 9052
rect 27274 9010 27318 9052
rect 27442 9010 27489 9052
rect 39103 9092 39150 9134
rect 39274 9092 39318 9134
rect 39442 9092 39489 9134
rect 39103 9052 39112 9092
rect 39274 9052 39276 9092
rect 39316 9052 39318 9092
rect 39480 9052 39489 9092
rect 39103 9010 39150 9052
rect 39274 9010 39318 9052
rect 39442 9010 39489 9052
rect 51103 9092 51150 9134
rect 51274 9092 51318 9134
rect 51442 9092 51489 9134
rect 51103 9052 51112 9092
rect 51274 9052 51276 9092
rect 51316 9052 51318 9092
rect 51480 9052 51489 9092
rect 51103 9010 51150 9052
rect 51274 9010 51318 9052
rect 51442 9010 51489 9052
rect 63103 9092 63150 9134
rect 63274 9092 63318 9134
rect 63442 9092 63489 9134
rect 63103 9052 63112 9092
rect 63274 9052 63276 9092
rect 63316 9052 63318 9092
rect 63480 9052 63489 9092
rect 63103 9010 63150 9052
rect 63274 9010 63318 9052
rect 63442 9010 63489 9052
rect 75103 9092 75150 9134
rect 75274 9092 75318 9134
rect 75442 9092 75489 9134
rect 75103 9052 75112 9092
rect 75274 9052 75276 9092
rect 75316 9052 75318 9092
rect 75480 9052 75489 9092
rect 75103 9010 75150 9052
rect 75274 9010 75318 9052
rect 75442 9010 75489 9052
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 16343 8336 16390 8378
rect 16514 8336 16558 8378
rect 16682 8336 16729 8378
rect 16343 8296 16352 8336
rect 16514 8296 16516 8336
rect 16556 8296 16558 8336
rect 16720 8296 16729 8336
rect 16343 8254 16390 8296
rect 16514 8254 16558 8296
rect 16682 8254 16729 8296
rect 28343 8336 28390 8378
rect 28514 8336 28558 8378
rect 28682 8336 28729 8378
rect 28343 8296 28352 8336
rect 28514 8296 28516 8336
rect 28556 8296 28558 8336
rect 28720 8296 28729 8336
rect 28343 8254 28390 8296
rect 28514 8254 28558 8296
rect 28682 8254 28729 8296
rect 40343 8336 40390 8378
rect 40514 8336 40558 8378
rect 40682 8336 40729 8378
rect 40343 8296 40352 8336
rect 40514 8296 40516 8336
rect 40556 8296 40558 8336
rect 40720 8296 40729 8336
rect 40343 8254 40390 8296
rect 40514 8254 40558 8296
rect 40682 8254 40729 8296
rect 52343 8336 52390 8378
rect 52514 8336 52558 8378
rect 52682 8336 52729 8378
rect 52343 8296 52352 8336
rect 52514 8296 52516 8336
rect 52556 8296 52558 8336
rect 52720 8296 52729 8336
rect 52343 8254 52390 8296
rect 52514 8254 52558 8296
rect 52682 8254 52729 8296
rect 64343 8336 64390 8378
rect 64514 8336 64558 8378
rect 64682 8336 64729 8378
rect 64343 8296 64352 8336
rect 64514 8296 64516 8336
rect 64556 8296 64558 8336
rect 64720 8296 64729 8336
rect 64343 8254 64390 8296
rect 64514 8254 64558 8296
rect 64682 8254 64729 8296
rect 76343 8336 76390 8378
rect 76514 8336 76558 8378
rect 76682 8336 76729 8378
rect 76343 8296 76352 8336
rect 76514 8296 76516 8336
rect 76556 8296 76558 8336
rect 76720 8296 76729 8336
rect 76343 8254 76390 8296
rect 76514 8254 76558 8296
rect 76682 8254 76729 8296
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 15103 7580 15150 7622
rect 15274 7580 15318 7622
rect 15442 7580 15489 7622
rect 15103 7540 15112 7580
rect 15274 7540 15276 7580
rect 15316 7540 15318 7580
rect 15480 7540 15489 7580
rect 15103 7498 15150 7540
rect 15274 7498 15318 7540
rect 15442 7498 15489 7540
rect 27103 7580 27150 7622
rect 27274 7580 27318 7622
rect 27442 7580 27489 7622
rect 27103 7540 27112 7580
rect 27274 7540 27276 7580
rect 27316 7540 27318 7580
rect 27480 7540 27489 7580
rect 27103 7498 27150 7540
rect 27274 7498 27318 7540
rect 27442 7498 27489 7540
rect 39103 7580 39150 7622
rect 39274 7580 39318 7622
rect 39442 7580 39489 7622
rect 39103 7540 39112 7580
rect 39274 7540 39276 7580
rect 39316 7540 39318 7580
rect 39480 7540 39489 7580
rect 39103 7498 39150 7540
rect 39274 7498 39318 7540
rect 39442 7498 39489 7540
rect 51103 7580 51150 7622
rect 51274 7580 51318 7622
rect 51442 7580 51489 7622
rect 51103 7540 51112 7580
rect 51274 7540 51276 7580
rect 51316 7540 51318 7580
rect 51480 7540 51489 7580
rect 51103 7498 51150 7540
rect 51274 7498 51318 7540
rect 51442 7498 51489 7540
rect 63103 7580 63150 7622
rect 63274 7580 63318 7622
rect 63442 7580 63489 7622
rect 63103 7540 63112 7580
rect 63274 7540 63276 7580
rect 63316 7540 63318 7580
rect 63480 7540 63489 7580
rect 63103 7498 63150 7540
rect 63274 7498 63318 7540
rect 63442 7498 63489 7540
rect 75103 7580 75150 7622
rect 75274 7580 75318 7622
rect 75442 7580 75489 7622
rect 75103 7540 75112 7580
rect 75274 7540 75276 7580
rect 75316 7540 75318 7580
rect 75480 7540 75489 7580
rect 75103 7498 75150 7540
rect 75274 7498 75318 7540
rect 75442 7498 75489 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 16343 6824 16390 6866
rect 16514 6824 16558 6866
rect 16682 6824 16729 6866
rect 16343 6784 16352 6824
rect 16514 6784 16516 6824
rect 16556 6784 16558 6824
rect 16720 6784 16729 6824
rect 16343 6742 16390 6784
rect 16514 6742 16558 6784
rect 16682 6742 16729 6784
rect 28343 6824 28390 6866
rect 28514 6824 28558 6866
rect 28682 6824 28729 6866
rect 28343 6784 28352 6824
rect 28514 6784 28516 6824
rect 28556 6784 28558 6824
rect 28720 6784 28729 6824
rect 28343 6742 28390 6784
rect 28514 6742 28558 6784
rect 28682 6742 28729 6784
rect 40343 6824 40390 6866
rect 40514 6824 40558 6866
rect 40682 6824 40729 6866
rect 40343 6784 40352 6824
rect 40514 6784 40516 6824
rect 40556 6784 40558 6824
rect 40720 6784 40729 6824
rect 40343 6742 40390 6784
rect 40514 6742 40558 6784
rect 40682 6742 40729 6784
rect 52343 6824 52390 6866
rect 52514 6824 52558 6866
rect 52682 6824 52729 6866
rect 52343 6784 52352 6824
rect 52514 6784 52516 6824
rect 52556 6784 52558 6824
rect 52720 6784 52729 6824
rect 52343 6742 52390 6784
rect 52514 6742 52558 6784
rect 52682 6742 52729 6784
rect 64343 6824 64390 6866
rect 64514 6824 64558 6866
rect 64682 6824 64729 6866
rect 64343 6784 64352 6824
rect 64514 6784 64516 6824
rect 64556 6784 64558 6824
rect 64720 6784 64729 6824
rect 64343 6742 64390 6784
rect 64514 6742 64558 6784
rect 64682 6742 64729 6784
rect 76343 6824 76390 6866
rect 76514 6824 76558 6866
rect 76682 6824 76729 6866
rect 76343 6784 76352 6824
rect 76514 6784 76516 6824
rect 76556 6784 76558 6824
rect 76720 6784 76729 6824
rect 76343 6742 76390 6784
rect 76514 6742 76558 6784
rect 76682 6742 76729 6784
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 15103 6068 15150 6110
rect 15274 6068 15318 6110
rect 15442 6068 15489 6110
rect 15103 6028 15112 6068
rect 15274 6028 15276 6068
rect 15316 6028 15318 6068
rect 15480 6028 15489 6068
rect 15103 5986 15150 6028
rect 15274 5986 15318 6028
rect 15442 5986 15489 6028
rect 27103 6068 27150 6110
rect 27274 6068 27318 6110
rect 27442 6068 27489 6110
rect 27103 6028 27112 6068
rect 27274 6028 27276 6068
rect 27316 6028 27318 6068
rect 27480 6028 27489 6068
rect 27103 5986 27150 6028
rect 27274 5986 27318 6028
rect 27442 5986 27489 6028
rect 39103 6068 39150 6110
rect 39274 6068 39318 6110
rect 39442 6068 39489 6110
rect 39103 6028 39112 6068
rect 39274 6028 39276 6068
rect 39316 6028 39318 6068
rect 39480 6028 39489 6068
rect 39103 5986 39150 6028
rect 39274 5986 39318 6028
rect 39442 5986 39489 6028
rect 51103 6068 51150 6110
rect 51274 6068 51318 6110
rect 51442 6068 51489 6110
rect 51103 6028 51112 6068
rect 51274 6028 51276 6068
rect 51316 6028 51318 6068
rect 51480 6028 51489 6068
rect 51103 5986 51150 6028
rect 51274 5986 51318 6028
rect 51442 5986 51489 6028
rect 63103 6068 63150 6110
rect 63274 6068 63318 6110
rect 63442 6068 63489 6110
rect 63103 6028 63112 6068
rect 63274 6028 63276 6068
rect 63316 6028 63318 6068
rect 63480 6028 63489 6068
rect 63103 5986 63150 6028
rect 63274 5986 63318 6028
rect 63442 5986 63489 6028
rect 75103 6068 75150 6110
rect 75274 6068 75318 6110
rect 75442 6068 75489 6110
rect 75103 6028 75112 6068
rect 75274 6028 75276 6068
rect 75316 6028 75318 6068
rect 75480 6028 75489 6068
rect 75103 5986 75150 6028
rect 75274 5986 75318 6028
rect 75442 5986 75489 6028
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 16343 5312 16390 5354
rect 16514 5312 16558 5354
rect 16682 5312 16729 5354
rect 16343 5272 16352 5312
rect 16514 5272 16516 5312
rect 16556 5272 16558 5312
rect 16720 5272 16729 5312
rect 16343 5230 16390 5272
rect 16514 5230 16558 5272
rect 16682 5230 16729 5272
rect 28343 5312 28390 5354
rect 28514 5312 28558 5354
rect 28682 5312 28729 5354
rect 28343 5272 28352 5312
rect 28514 5272 28516 5312
rect 28556 5272 28558 5312
rect 28720 5272 28729 5312
rect 28343 5230 28390 5272
rect 28514 5230 28558 5272
rect 28682 5230 28729 5272
rect 40343 5312 40390 5354
rect 40514 5312 40558 5354
rect 40682 5312 40729 5354
rect 40343 5272 40352 5312
rect 40514 5272 40516 5312
rect 40556 5272 40558 5312
rect 40720 5272 40729 5312
rect 40343 5230 40390 5272
rect 40514 5230 40558 5272
rect 40682 5230 40729 5272
rect 52343 5312 52390 5354
rect 52514 5312 52558 5354
rect 52682 5312 52729 5354
rect 52343 5272 52352 5312
rect 52514 5272 52516 5312
rect 52556 5272 52558 5312
rect 52720 5272 52729 5312
rect 52343 5230 52390 5272
rect 52514 5230 52558 5272
rect 52682 5230 52729 5272
rect 64343 5312 64390 5354
rect 64514 5312 64558 5354
rect 64682 5312 64729 5354
rect 64343 5272 64352 5312
rect 64514 5272 64516 5312
rect 64556 5272 64558 5312
rect 64720 5272 64729 5312
rect 64343 5230 64390 5272
rect 64514 5230 64558 5272
rect 64682 5230 64729 5272
rect 76343 5312 76390 5354
rect 76514 5312 76558 5354
rect 76682 5312 76729 5354
rect 76343 5272 76352 5312
rect 76514 5272 76516 5312
rect 76556 5272 76558 5312
rect 76720 5272 76729 5312
rect 76343 5230 76390 5272
rect 76514 5230 76558 5272
rect 76682 5230 76729 5272
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 15103 4556 15150 4598
rect 15274 4556 15318 4598
rect 15442 4556 15489 4598
rect 15103 4516 15112 4556
rect 15274 4516 15276 4556
rect 15316 4516 15318 4556
rect 15480 4516 15489 4556
rect 15103 4474 15150 4516
rect 15274 4474 15318 4516
rect 15442 4474 15489 4516
rect 27103 4556 27150 4598
rect 27274 4556 27318 4598
rect 27442 4556 27489 4598
rect 27103 4516 27112 4556
rect 27274 4516 27276 4556
rect 27316 4516 27318 4556
rect 27480 4516 27489 4556
rect 27103 4474 27150 4516
rect 27274 4474 27318 4516
rect 27442 4474 27489 4516
rect 39103 4556 39150 4598
rect 39274 4556 39318 4598
rect 39442 4556 39489 4598
rect 39103 4516 39112 4556
rect 39274 4516 39276 4556
rect 39316 4516 39318 4556
rect 39480 4516 39489 4556
rect 39103 4474 39150 4516
rect 39274 4474 39318 4516
rect 39442 4474 39489 4516
rect 51103 4556 51150 4598
rect 51274 4556 51318 4598
rect 51442 4556 51489 4598
rect 51103 4516 51112 4556
rect 51274 4516 51276 4556
rect 51316 4516 51318 4556
rect 51480 4516 51489 4556
rect 51103 4474 51150 4516
rect 51274 4474 51318 4516
rect 51442 4474 51489 4516
rect 63103 4556 63150 4598
rect 63274 4556 63318 4598
rect 63442 4556 63489 4598
rect 63103 4516 63112 4556
rect 63274 4516 63276 4556
rect 63316 4516 63318 4556
rect 63480 4516 63489 4556
rect 63103 4474 63150 4516
rect 63274 4474 63318 4516
rect 63442 4474 63489 4516
rect 75103 4556 75150 4598
rect 75274 4556 75318 4598
rect 75442 4556 75489 4598
rect 75103 4516 75112 4556
rect 75274 4516 75276 4556
rect 75316 4516 75318 4556
rect 75480 4516 75489 4556
rect 75103 4474 75150 4516
rect 75274 4474 75318 4516
rect 75442 4474 75489 4516
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 16343 3800 16390 3842
rect 16514 3800 16558 3842
rect 16682 3800 16729 3842
rect 16343 3760 16352 3800
rect 16514 3760 16516 3800
rect 16556 3760 16558 3800
rect 16720 3760 16729 3800
rect 16343 3718 16390 3760
rect 16514 3718 16558 3760
rect 16682 3718 16729 3760
rect 28343 3800 28390 3842
rect 28514 3800 28558 3842
rect 28682 3800 28729 3842
rect 28343 3760 28352 3800
rect 28514 3760 28516 3800
rect 28556 3760 28558 3800
rect 28720 3760 28729 3800
rect 28343 3718 28390 3760
rect 28514 3718 28558 3760
rect 28682 3718 28729 3760
rect 40343 3800 40390 3842
rect 40514 3800 40558 3842
rect 40682 3800 40729 3842
rect 40343 3760 40352 3800
rect 40514 3760 40516 3800
rect 40556 3760 40558 3800
rect 40720 3760 40729 3800
rect 40343 3718 40390 3760
rect 40514 3718 40558 3760
rect 40682 3718 40729 3760
rect 52343 3800 52390 3842
rect 52514 3800 52558 3842
rect 52682 3800 52729 3842
rect 52343 3760 52352 3800
rect 52514 3760 52516 3800
rect 52556 3760 52558 3800
rect 52720 3760 52729 3800
rect 52343 3718 52390 3760
rect 52514 3718 52558 3760
rect 52682 3718 52729 3760
rect 64343 3800 64390 3842
rect 64514 3800 64558 3842
rect 64682 3800 64729 3842
rect 64343 3760 64352 3800
rect 64514 3760 64516 3800
rect 64556 3760 64558 3800
rect 64720 3760 64729 3800
rect 64343 3718 64390 3760
rect 64514 3718 64558 3760
rect 64682 3718 64729 3760
rect 76343 3800 76390 3842
rect 76514 3800 76558 3842
rect 76682 3800 76729 3842
rect 76343 3760 76352 3800
rect 76514 3760 76516 3800
rect 76556 3760 76558 3800
rect 76720 3760 76729 3800
rect 76343 3718 76390 3760
rect 76514 3718 76558 3760
rect 76682 3718 76729 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 15103 3044 15150 3086
rect 15274 3044 15318 3086
rect 15442 3044 15489 3086
rect 15103 3004 15112 3044
rect 15274 3004 15276 3044
rect 15316 3004 15318 3044
rect 15480 3004 15489 3044
rect 15103 2962 15150 3004
rect 15274 2962 15318 3004
rect 15442 2962 15489 3004
rect 27103 3044 27150 3086
rect 27274 3044 27318 3086
rect 27442 3044 27489 3086
rect 27103 3004 27112 3044
rect 27274 3004 27276 3044
rect 27316 3004 27318 3044
rect 27480 3004 27489 3044
rect 27103 2962 27150 3004
rect 27274 2962 27318 3004
rect 27442 2962 27489 3004
rect 39103 3044 39150 3086
rect 39274 3044 39318 3086
rect 39442 3044 39489 3086
rect 39103 3004 39112 3044
rect 39274 3004 39276 3044
rect 39316 3004 39318 3044
rect 39480 3004 39489 3044
rect 39103 2962 39150 3004
rect 39274 2962 39318 3004
rect 39442 2962 39489 3004
rect 51103 3044 51150 3086
rect 51274 3044 51318 3086
rect 51442 3044 51489 3086
rect 51103 3004 51112 3044
rect 51274 3004 51276 3044
rect 51316 3004 51318 3044
rect 51480 3004 51489 3044
rect 51103 2962 51150 3004
rect 51274 2962 51318 3004
rect 51442 2962 51489 3004
rect 63103 3044 63150 3086
rect 63274 3044 63318 3086
rect 63442 3044 63489 3086
rect 63103 3004 63112 3044
rect 63274 3004 63276 3044
rect 63316 3004 63318 3044
rect 63480 3004 63489 3044
rect 63103 2962 63150 3004
rect 63274 2962 63318 3004
rect 63442 2962 63489 3004
rect 75103 3044 75150 3086
rect 75274 3044 75318 3086
rect 75442 3044 75489 3086
rect 75103 3004 75112 3044
rect 75274 3004 75276 3044
rect 75316 3004 75318 3044
rect 75480 3004 75489 3044
rect 75103 2962 75150 3004
rect 75274 2962 75318 3004
rect 75442 2962 75489 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 16343 2288 16390 2330
rect 16514 2288 16558 2330
rect 16682 2288 16729 2330
rect 16343 2248 16352 2288
rect 16514 2248 16516 2288
rect 16556 2248 16558 2288
rect 16720 2248 16729 2288
rect 16343 2206 16390 2248
rect 16514 2206 16558 2248
rect 16682 2206 16729 2248
rect 28343 2288 28390 2330
rect 28514 2288 28558 2330
rect 28682 2288 28729 2330
rect 28343 2248 28352 2288
rect 28514 2248 28516 2288
rect 28556 2248 28558 2288
rect 28720 2248 28729 2288
rect 28343 2206 28390 2248
rect 28514 2206 28558 2248
rect 28682 2206 28729 2248
rect 40343 2288 40390 2330
rect 40514 2288 40558 2330
rect 40682 2288 40729 2330
rect 40343 2248 40352 2288
rect 40514 2248 40516 2288
rect 40556 2248 40558 2288
rect 40720 2248 40729 2288
rect 40343 2206 40390 2248
rect 40514 2206 40558 2248
rect 40682 2206 40729 2248
rect 52343 2288 52390 2330
rect 52514 2288 52558 2330
rect 52682 2288 52729 2330
rect 52343 2248 52352 2288
rect 52514 2248 52516 2288
rect 52556 2248 52558 2288
rect 52720 2248 52729 2288
rect 52343 2206 52390 2248
rect 52514 2206 52558 2248
rect 52682 2206 52729 2248
rect 64343 2288 64390 2330
rect 64514 2288 64558 2330
rect 64682 2288 64729 2330
rect 64343 2248 64352 2288
rect 64514 2248 64516 2288
rect 64556 2248 64558 2288
rect 64720 2248 64729 2288
rect 64343 2206 64390 2248
rect 64514 2206 64558 2248
rect 64682 2206 64729 2248
rect 76343 2288 76390 2330
rect 76514 2288 76558 2330
rect 76682 2288 76729 2330
rect 76343 2248 76352 2288
rect 76514 2248 76516 2288
rect 76556 2248 76558 2288
rect 76720 2248 76729 2288
rect 76343 2206 76390 2248
rect 76514 2206 76558 2248
rect 76682 2206 76729 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 15103 1532 15150 1574
rect 15274 1532 15318 1574
rect 15442 1532 15489 1574
rect 15103 1492 15112 1532
rect 15274 1492 15276 1532
rect 15316 1492 15318 1532
rect 15480 1492 15489 1532
rect 15103 1450 15150 1492
rect 15274 1450 15318 1492
rect 15442 1450 15489 1492
rect 27103 1532 27150 1574
rect 27274 1532 27318 1574
rect 27442 1532 27489 1574
rect 27103 1492 27112 1532
rect 27274 1492 27276 1532
rect 27316 1492 27318 1532
rect 27480 1492 27489 1532
rect 27103 1450 27150 1492
rect 27274 1450 27318 1492
rect 27442 1450 27489 1492
rect 39103 1532 39150 1574
rect 39274 1532 39318 1574
rect 39442 1532 39489 1574
rect 39103 1492 39112 1532
rect 39274 1492 39276 1532
rect 39316 1492 39318 1532
rect 39480 1492 39489 1532
rect 39103 1450 39150 1492
rect 39274 1450 39318 1492
rect 39442 1450 39489 1492
rect 51103 1532 51150 1574
rect 51274 1532 51318 1574
rect 51442 1532 51489 1574
rect 51103 1492 51112 1532
rect 51274 1492 51276 1532
rect 51316 1492 51318 1532
rect 51480 1492 51489 1532
rect 51103 1450 51150 1492
rect 51274 1450 51318 1492
rect 51442 1450 51489 1492
rect 63103 1532 63150 1574
rect 63274 1532 63318 1574
rect 63442 1532 63489 1574
rect 63103 1492 63112 1532
rect 63274 1492 63276 1532
rect 63316 1492 63318 1532
rect 63480 1492 63489 1532
rect 63103 1450 63150 1492
rect 63274 1450 63318 1492
rect 63442 1450 63489 1492
rect 75103 1532 75150 1574
rect 75274 1532 75318 1574
rect 75442 1532 75489 1574
rect 75103 1492 75112 1532
rect 75274 1492 75276 1532
rect 75316 1492 75318 1532
rect 75480 1492 75489 1532
rect 75103 1450 75150 1492
rect 75274 1450 75318 1492
rect 75442 1450 75489 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 16343 776 16390 818
rect 16514 776 16558 818
rect 16682 776 16729 818
rect 16343 736 16352 776
rect 16514 736 16516 776
rect 16556 736 16558 776
rect 16720 736 16729 776
rect 16343 694 16390 736
rect 16514 694 16558 736
rect 16682 694 16729 736
rect 28343 776 28390 818
rect 28514 776 28558 818
rect 28682 776 28729 818
rect 28343 736 28352 776
rect 28514 736 28516 776
rect 28556 736 28558 776
rect 28720 736 28729 776
rect 28343 694 28390 736
rect 28514 694 28558 736
rect 28682 694 28729 736
rect 40343 776 40390 818
rect 40514 776 40558 818
rect 40682 776 40729 818
rect 40343 736 40352 776
rect 40514 736 40516 776
rect 40556 736 40558 776
rect 40720 736 40729 776
rect 40343 694 40390 736
rect 40514 694 40558 736
rect 40682 694 40729 736
rect 52343 776 52390 818
rect 52514 776 52558 818
rect 52682 776 52729 818
rect 52343 736 52352 776
rect 52514 736 52516 776
rect 52556 736 52558 776
rect 52720 736 52729 776
rect 52343 694 52390 736
rect 52514 694 52558 736
rect 52682 694 52729 736
rect 64343 776 64390 818
rect 64514 776 64558 818
rect 64682 776 64729 818
rect 64343 736 64352 776
rect 64514 736 64516 776
rect 64556 736 64558 776
rect 64720 736 64729 776
rect 64343 694 64390 736
rect 64514 694 64558 736
rect 64682 694 64729 736
rect 76343 776 76390 818
rect 76514 776 76558 818
rect 76682 776 76729 818
rect 76343 736 76352 776
rect 76514 736 76516 776
rect 76556 736 76558 776
rect 76720 736 76729 776
rect 76343 694 76390 736
rect 76514 694 76558 736
rect 76682 694 76729 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 16390 38576 16514 38618
rect 16558 38576 16682 38618
rect 16390 38536 16392 38576
rect 16392 38536 16434 38576
rect 16434 38536 16474 38576
rect 16474 38536 16514 38576
rect 16558 38536 16598 38576
rect 16598 38536 16638 38576
rect 16638 38536 16680 38576
rect 16680 38536 16682 38576
rect 16390 38494 16514 38536
rect 16558 38494 16682 38536
rect 28390 38576 28514 38618
rect 28558 38576 28682 38618
rect 28390 38536 28392 38576
rect 28392 38536 28434 38576
rect 28434 38536 28474 38576
rect 28474 38536 28514 38576
rect 28558 38536 28598 38576
rect 28598 38536 28638 38576
rect 28638 38536 28680 38576
rect 28680 38536 28682 38576
rect 28390 38494 28514 38536
rect 28558 38494 28682 38536
rect 40390 38576 40514 38618
rect 40558 38576 40682 38618
rect 40390 38536 40392 38576
rect 40392 38536 40434 38576
rect 40434 38536 40474 38576
rect 40474 38536 40514 38576
rect 40558 38536 40598 38576
rect 40598 38536 40638 38576
rect 40638 38536 40680 38576
rect 40680 38536 40682 38576
rect 40390 38494 40514 38536
rect 40558 38494 40682 38536
rect 52390 38576 52514 38618
rect 52558 38576 52682 38618
rect 52390 38536 52392 38576
rect 52392 38536 52434 38576
rect 52434 38536 52474 38576
rect 52474 38536 52514 38576
rect 52558 38536 52598 38576
rect 52598 38536 52638 38576
rect 52638 38536 52680 38576
rect 52680 38536 52682 38576
rect 52390 38494 52514 38536
rect 52558 38494 52682 38536
rect 64390 38576 64514 38618
rect 64558 38576 64682 38618
rect 64390 38536 64392 38576
rect 64392 38536 64434 38576
rect 64434 38536 64474 38576
rect 64474 38536 64514 38576
rect 64558 38536 64598 38576
rect 64598 38536 64638 38576
rect 64638 38536 64680 38576
rect 64680 38536 64682 38576
rect 64390 38494 64514 38536
rect 64558 38494 64682 38536
rect 76390 38576 76514 38618
rect 76558 38576 76682 38618
rect 76390 38536 76392 38576
rect 76392 38536 76434 38576
rect 76434 38536 76474 38576
rect 76474 38536 76514 38576
rect 76558 38536 76598 38576
rect 76598 38536 76638 38576
rect 76638 38536 76680 38576
rect 76680 38536 76682 38576
rect 76390 38494 76514 38536
rect 76558 38494 76682 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 15150 37820 15274 37862
rect 15318 37820 15442 37862
rect 15150 37780 15152 37820
rect 15152 37780 15194 37820
rect 15194 37780 15234 37820
rect 15234 37780 15274 37820
rect 15318 37780 15358 37820
rect 15358 37780 15398 37820
rect 15398 37780 15440 37820
rect 15440 37780 15442 37820
rect 15150 37738 15274 37780
rect 15318 37738 15442 37780
rect 27150 37820 27274 37862
rect 27318 37820 27442 37862
rect 27150 37780 27152 37820
rect 27152 37780 27194 37820
rect 27194 37780 27234 37820
rect 27234 37780 27274 37820
rect 27318 37780 27358 37820
rect 27358 37780 27398 37820
rect 27398 37780 27440 37820
rect 27440 37780 27442 37820
rect 27150 37738 27274 37780
rect 27318 37738 27442 37780
rect 39150 37820 39274 37862
rect 39318 37820 39442 37862
rect 39150 37780 39152 37820
rect 39152 37780 39194 37820
rect 39194 37780 39234 37820
rect 39234 37780 39274 37820
rect 39318 37780 39358 37820
rect 39358 37780 39398 37820
rect 39398 37780 39440 37820
rect 39440 37780 39442 37820
rect 39150 37738 39274 37780
rect 39318 37738 39442 37780
rect 51150 37820 51274 37862
rect 51318 37820 51442 37862
rect 51150 37780 51152 37820
rect 51152 37780 51194 37820
rect 51194 37780 51234 37820
rect 51234 37780 51274 37820
rect 51318 37780 51358 37820
rect 51358 37780 51398 37820
rect 51398 37780 51440 37820
rect 51440 37780 51442 37820
rect 51150 37738 51274 37780
rect 51318 37738 51442 37780
rect 63150 37820 63274 37862
rect 63318 37820 63442 37862
rect 63150 37780 63152 37820
rect 63152 37780 63194 37820
rect 63194 37780 63234 37820
rect 63234 37780 63274 37820
rect 63318 37780 63358 37820
rect 63358 37780 63398 37820
rect 63398 37780 63440 37820
rect 63440 37780 63442 37820
rect 63150 37738 63274 37780
rect 63318 37738 63442 37780
rect 75150 37820 75274 37862
rect 75318 37820 75442 37862
rect 75150 37780 75152 37820
rect 75152 37780 75194 37820
rect 75194 37780 75234 37820
rect 75234 37780 75274 37820
rect 75318 37780 75358 37820
rect 75358 37780 75398 37820
rect 75398 37780 75440 37820
rect 75440 37780 75442 37820
rect 75150 37738 75274 37780
rect 75318 37738 75442 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 16390 37064 16514 37106
rect 16558 37064 16682 37106
rect 16390 37024 16392 37064
rect 16392 37024 16434 37064
rect 16434 37024 16474 37064
rect 16474 37024 16514 37064
rect 16558 37024 16598 37064
rect 16598 37024 16638 37064
rect 16638 37024 16680 37064
rect 16680 37024 16682 37064
rect 16390 36982 16514 37024
rect 16558 36982 16682 37024
rect 28390 37064 28514 37106
rect 28558 37064 28682 37106
rect 28390 37024 28392 37064
rect 28392 37024 28434 37064
rect 28434 37024 28474 37064
rect 28474 37024 28514 37064
rect 28558 37024 28598 37064
rect 28598 37024 28638 37064
rect 28638 37024 28680 37064
rect 28680 37024 28682 37064
rect 28390 36982 28514 37024
rect 28558 36982 28682 37024
rect 40390 37064 40514 37106
rect 40558 37064 40682 37106
rect 40390 37024 40392 37064
rect 40392 37024 40434 37064
rect 40434 37024 40474 37064
rect 40474 37024 40514 37064
rect 40558 37024 40598 37064
rect 40598 37024 40638 37064
rect 40638 37024 40680 37064
rect 40680 37024 40682 37064
rect 40390 36982 40514 37024
rect 40558 36982 40682 37024
rect 52390 37064 52514 37106
rect 52558 37064 52682 37106
rect 52390 37024 52392 37064
rect 52392 37024 52434 37064
rect 52434 37024 52474 37064
rect 52474 37024 52514 37064
rect 52558 37024 52598 37064
rect 52598 37024 52638 37064
rect 52638 37024 52680 37064
rect 52680 37024 52682 37064
rect 52390 36982 52514 37024
rect 52558 36982 52682 37024
rect 64390 37064 64514 37106
rect 64558 37064 64682 37106
rect 64390 37024 64392 37064
rect 64392 37024 64434 37064
rect 64434 37024 64474 37064
rect 64474 37024 64514 37064
rect 64558 37024 64598 37064
rect 64598 37024 64638 37064
rect 64638 37024 64680 37064
rect 64680 37024 64682 37064
rect 64390 36982 64514 37024
rect 64558 36982 64682 37024
rect 76390 37064 76514 37106
rect 76558 37064 76682 37106
rect 76390 37024 76392 37064
rect 76392 37024 76434 37064
rect 76434 37024 76474 37064
rect 76474 37024 76514 37064
rect 76558 37024 76598 37064
rect 76598 37024 76638 37064
rect 76638 37024 76680 37064
rect 76680 37024 76682 37064
rect 76390 36982 76514 37024
rect 76558 36982 76682 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 15150 36308 15274 36350
rect 15318 36308 15442 36350
rect 15150 36268 15152 36308
rect 15152 36268 15194 36308
rect 15194 36268 15234 36308
rect 15234 36268 15274 36308
rect 15318 36268 15358 36308
rect 15358 36268 15398 36308
rect 15398 36268 15440 36308
rect 15440 36268 15442 36308
rect 15150 36226 15274 36268
rect 15318 36226 15442 36268
rect 27150 36308 27274 36350
rect 27318 36308 27442 36350
rect 27150 36268 27152 36308
rect 27152 36268 27194 36308
rect 27194 36268 27234 36308
rect 27234 36268 27274 36308
rect 27318 36268 27358 36308
rect 27358 36268 27398 36308
rect 27398 36268 27440 36308
rect 27440 36268 27442 36308
rect 27150 36226 27274 36268
rect 27318 36226 27442 36268
rect 39150 36308 39274 36350
rect 39318 36308 39442 36350
rect 39150 36268 39152 36308
rect 39152 36268 39194 36308
rect 39194 36268 39234 36308
rect 39234 36268 39274 36308
rect 39318 36268 39358 36308
rect 39358 36268 39398 36308
rect 39398 36268 39440 36308
rect 39440 36268 39442 36308
rect 39150 36226 39274 36268
rect 39318 36226 39442 36268
rect 51150 36308 51274 36350
rect 51318 36308 51442 36350
rect 51150 36268 51152 36308
rect 51152 36268 51194 36308
rect 51194 36268 51234 36308
rect 51234 36268 51274 36308
rect 51318 36268 51358 36308
rect 51358 36268 51398 36308
rect 51398 36268 51440 36308
rect 51440 36268 51442 36308
rect 51150 36226 51274 36268
rect 51318 36226 51442 36268
rect 63150 36308 63274 36350
rect 63318 36308 63442 36350
rect 63150 36268 63152 36308
rect 63152 36268 63194 36308
rect 63194 36268 63234 36308
rect 63234 36268 63274 36308
rect 63318 36268 63358 36308
rect 63358 36268 63398 36308
rect 63398 36268 63440 36308
rect 63440 36268 63442 36308
rect 63150 36226 63274 36268
rect 63318 36226 63442 36268
rect 75150 36308 75274 36350
rect 75318 36308 75442 36350
rect 75150 36268 75152 36308
rect 75152 36268 75194 36308
rect 75194 36268 75234 36308
rect 75234 36268 75274 36308
rect 75318 36268 75358 36308
rect 75358 36268 75398 36308
rect 75398 36268 75440 36308
rect 75440 36268 75442 36308
rect 75150 36226 75274 36268
rect 75318 36226 75442 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 16390 35552 16514 35594
rect 16558 35552 16682 35594
rect 16390 35512 16392 35552
rect 16392 35512 16434 35552
rect 16434 35512 16474 35552
rect 16474 35512 16514 35552
rect 16558 35512 16598 35552
rect 16598 35512 16638 35552
rect 16638 35512 16680 35552
rect 16680 35512 16682 35552
rect 16390 35470 16514 35512
rect 16558 35470 16682 35512
rect 28390 35552 28514 35594
rect 28558 35552 28682 35594
rect 28390 35512 28392 35552
rect 28392 35512 28434 35552
rect 28434 35512 28474 35552
rect 28474 35512 28514 35552
rect 28558 35512 28598 35552
rect 28598 35512 28638 35552
rect 28638 35512 28680 35552
rect 28680 35512 28682 35552
rect 28390 35470 28514 35512
rect 28558 35470 28682 35512
rect 40390 35552 40514 35594
rect 40558 35552 40682 35594
rect 40390 35512 40392 35552
rect 40392 35512 40434 35552
rect 40434 35512 40474 35552
rect 40474 35512 40514 35552
rect 40558 35512 40598 35552
rect 40598 35512 40638 35552
rect 40638 35512 40680 35552
rect 40680 35512 40682 35552
rect 40390 35470 40514 35512
rect 40558 35470 40682 35512
rect 52390 35552 52514 35594
rect 52558 35552 52682 35594
rect 52390 35512 52392 35552
rect 52392 35512 52434 35552
rect 52434 35512 52474 35552
rect 52474 35512 52514 35552
rect 52558 35512 52598 35552
rect 52598 35512 52638 35552
rect 52638 35512 52680 35552
rect 52680 35512 52682 35552
rect 52390 35470 52514 35512
rect 52558 35470 52682 35512
rect 64390 35552 64514 35594
rect 64558 35552 64682 35594
rect 64390 35512 64392 35552
rect 64392 35512 64434 35552
rect 64434 35512 64474 35552
rect 64474 35512 64514 35552
rect 64558 35512 64598 35552
rect 64598 35512 64638 35552
rect 64638 35512 64680 35552
rect 64680 35512 64682 35552
rect 64390 35470 64514 35512
rect 64558 35470 64682 35512
rect 76390 35552 76514 35594
rect 76558 35552 76682 35594
rect 76390 35512 76392 35552
rect 76392 35512 76434 35552
rect 76434 35512 76474 35552
rect 76474 35512 76514 35552
rect 76558 35512 76598 35552
rect 76598 35512 76638 35552
rect 76638 35512 76680 35552
rect 76680 35512 76682 35552
rect 76390 35470 76514 35512
rect 76558 35470 76682 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 15150 34796 15274 34838
rect 15318 34796 15442 34838
rect 15150 34756 15152 34796
rect 15152 34756 15194 34796
rect 15194 34756 15234 34796
rect 15234 34756 15274 34796
rect 15318 34756 15358 34796
rect 15358 34756 15398 34796
rect 15398 34756 15440 34796
rect 15440 34756 15442 34796
rect 15150 34714 15274 34756
rect 15318 34714 15442 34756
rect 27150 34796 27274 34838
rect 27318 34796 27442 34838
rect 27150 34756 27152 34796
rect 27152 34756 27194 34796
rect 27194 34756 27234 34796
rect 27234 34756 27274 34796
rect 27318 34756 27358 34796
rect 27358 34756 27398 34796
rect 27398 34756 27440 34796
rect 27440 34756 27442 34796
rect 27150 34714 27274 34756
rect 27318 34714 27442 34756
rect 39150 34796 39274 34838
rect 39318 34796 39442 34838
rect 39150 34756 39152 34796
rect 39152 34756 39194 34796
rect 39194 34756 39234 34796
rect 39234 34756 39274 34796
rect 39318 34756 39358 34796
rect 39358 34756 39398 34796
rect 39398 34756 39440 34796
rect 39440 34756 39442 34796
rect 39150 34714 39274 34756
rect 39318 34714 39442 34756
rect 51150 34796 51274 34838
rect 51318 34796 51442 34838
rect 51150 34756 51152 34796
rect 51152 34756 51194 34796
rect 51194 34756 51234 34796
rect 51234 34756 51274 34796
rect 51318 34756 51358 34796
rect 51358 34756 51398 34796
rect 51398 34756 51440 34796
rect 51440 34756 51442 34796
rect 51150 34714 51274 34756
rect 51318 34714 51442 34756
rect 63150 34796 63274 34838
rect 63318 34796 63442 34838
rect 63150 34756 63152 34796
rect 63152 34756 63194 34796
rect 63194 34756 63234 34796
rect 63234 34756 63274 34796
rect 63318 34756 63358 34796
rect 63358 34756 63398 34796
rect 63398 34756 63440 34796
rect 63440 34756 63442 34796
rect 63150 34714 63274 34756
rect 63318 34714 63442 34756
rect 75150 34796 75274 34838
rect 75318 34796 75442 34838
rect 75150 34756 75152 34796
rect 75152 34756 75194 34796
rect 75194 34756 75234 34796
rect 75234 34756 75274 34796
rect 75318 34756 75358 34796
rect 75358 34756 75398 34796
rect 75398 34756 75440 34796
rect 75440 34756 75442 34796
rect 75150 34714 75274 34756
rect 75318 34714 75442 34756
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 16390 34040 16514 34082
rect 16558 34040 16682 34082
rect 16390 34000 16392 34040
rect 16392 34000 16434 34040
rect 16434 34000 16474 34040
rect 16474 34000 16514 34040
rect 16558 34000 16598 34040
rect 16598 34000 16638 34040
rect 16638 34000 16680 34040
rect 16680 34000 16682 34040
rect 16390 33958 16514 34000
rect 16558 33958 16682 34000
rect 28390 34040 28514 34082
rect 28558 34040 28682 34082
rect 28390 34000 28392 34040
rect 28392 34000 28434 34040
rect 28434 34000 28474 34040
rect 28474 34000 28514 34040
rect 28558 34000 28598 34040
rect 28598 34000 28638 34040
rect 28638 34000 28680 34040
rect 28680 34000 28682 34040
rect 28390 33958 28514 34000
rect 28558 33958 28682 34000
rect 40390 34040 40514 34082
rect 40558 34040 40682 34082
rect 40390 34000 40392 34040
rect 40392 34000 40434 34040
rect 40434 34000 40474 34040
rect 40474 34000 40514 34040
rect 40558 34000 40598 34040
rect 40598 34000 40638 34040
rect 40638 34000 40680 34040
rect 40680 34000 40682 34040
rect 40390 33958 40514 34000
rect 40558 33958 40682 34000
rect 52390 34040 52514 34082
rect 52558 34040 52682 34082
rect 52390 34000 52392 34040
rect 52392 34000 52434 34040
rect 52434 34000 52474 34040
rect 52474 34000 52514 34040
rect 52558 34000 52598 34040
rect 52598 34000 52638 34040
rect 52638 34000 52680 34040
rect 52680 34000 52682 34040
rect 52390 33958 52514 34000
rect 52558 33958 52682 34000
rect 64390 34040 64514 34082
rect 64558 34040 64682 34082
rect 64390 34000 64392 34040
rect 64392 34000 64434 34040
rect 64434 34000 64474 34040
rect 64474 34000 64514 34040
rect 64558 34000 64598 34040
rect 64598 34000 64638 34040
rect 64638 34000 64680 34040
rect 64680 34000 64682 34040
rect 64390 33958 64514 34000
rect 64558 33958 64682 34000
rect 76390 34040 76514 34082
rect 76558 34040 76682 34082
rect 76390 34000 76392 34040
rect 76392 34000 76434 34040
rect 76434 34000 76474 34040
rect 76474 34000 76514 34040
rect 76558 34000 76598 34040
rect 76598 34000 76638 34040
rect 76638 34000 76680 34040
rect 76680 34000 76682 34040
rect 76390 33958 76514 34000
rect 76558 33958 76682 34000
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 15150 33284 15274 33326
rect 15318 33284 15442 33326
rect 15150 33244 15152 33284
rect 15152 33244 15194 33284
rect 15194 33244 15234 33284
rect 15234 33244 15274 33284
rect 15318 33244 15358 33284
rect 15358 33244 15398 33284
rect 15398 33244 15440 33284
rect 15440 33244 15442 33284
rect 15150 33202 15274 33244
rect 15318 33202 15442 33244
rect 27150 33284 27274 33326
rect 27318 33284 27442 33326
rect 27150 33244 27152 33284
rect 27152 33244 27194 33284
rect 27194 33244 27234 33284
rect 27234 33244 27274 33284
rect 27318 33244 27358 33284
rect 27358 33244 27398 33284
rect 27398 33244 27440 33284
rect 27440 33244 27442 33284
rect 27150 33202 27274 33244
rect 27318 33202 27442 33244
rect 39150 33284 39274 33326
rect 39318 33284 39442 33326
rect 39150 33244 39152 33284
rect 39152 33244 39194 33284
rect 39194 33244 39234 33284
rect 39234 33244 39274 33284
rect 39318 33244 39358 33284
rect 39358 33244 39398 33284
rect 39398 33244 39440 33284
rect 39440 33244 39442 33284
rect 39150 33202 39274 33244
rect 39318 33202 39442 33244
rect 51150 33284 51274 33326
rect 51318 33284 51442 33326
rect 51150 33244 51152 33284
rect 51152 33244 51194 33284
rect 51194 33244 51234 33284
rect 51234 33244 51274 33284
rect 51318 33244 51358 33284
rect 51358 33244 51398 33284
rect 51398 33244 51440 33284
rect 51440 33244 51442 33284
rect 51150 33202 51274 33244
rect 51318 33202 51442 33244
rect 63150 33284 63274 33326
rect 63318 33284 63442 33326
rect 63150 33244 63152 33284
rect 63152 33244 63194 33284
rect 63194 33244 63234 33284
rect 63234 33244 63274 33284
rect 63318 33244 63358 33284
rect 63358 33244 63398 33284
rect 63398 33244 63440 33284
rect 63440 33244 63442 33284
rect 63150 33202 63274 33244
rect 63318 33202 63442 33244
rect 75150 33284 75274 33326
rect 75318 33284 75442 33326
rect 75150 33244 75152 33284
rect 75152 33244 75194 33284
rect 75194 33244 75234 33284
rect 75234 33244 75274 33284
rect 75318 33244 75358 33284
rect 75358 33244 75398 33284
rect 75398 33244 75440 33284
rect 75440 33244 75442 33284
rect 75150 33202 75274 33244
rect 75318 33202 75442 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 16390 32528 16514 32570
rect 16558 32528 16682 32570
rect 16390 32488 16392 32528
rect 16392 32488 16434 32528
rect 16434 32488 16474 32528
rect 16474 32488 16514 32528
rect 16558 32488 16598 32528
rect 16598 32488 16638 32528
rect 16638 32488 16680 32528
rect 16680 32488 16682 32528
rect 16390 32446 16514 32488
rect 16558 32446 16682 32488
rect 28390 32528 28514 32570
rect 28558 32528 28682 32570
rect 28390 32488 28392 32528
rect 28392 32488 28434 32528
rect 28434 32488 28474 32528
rect 28474 32488 28514 32528
rect 28558 32488 28598 32528
rect 28598 32488 28638 32528
rect 28638 32488 28680 32528
rect 28680 32488 28682 32528
rect 28390 32446 28514 32488
rect 28558 32446 28682 32488
rect 40390 32528 40514 32570
rect 40558 32528 40682 32570
rect 40390 32488 40392 32528
rect 40392 32488 40434 32528
rect 40434 32488 40474 32528
rect 40474 32488 40514 32528
rect 40558 32488 40598 32528
rect 40598 32488 40638 32528
rect 40638 32488 40680 32528
rect 40680 32488 40682 32528
rect 40390 32446 40514 32488
rect 40558 32446 40682 32488
rect 52390 32528 52514 32570
rect 52558 32528 52682 32570
rect 52390 32488 52392 32528
rect 52392 32488 52434 32528
rect 52434 32488 52474 32528
rect 52474 32488 52514 32528
rect 52558 32488 52598 32528
rect 52598 32488 52638 32528
rect 52638 32488 52680 32528
rect 52680 32488 52682 32528
rect 52390 32446 52514 32488
rect 52558 32446 52682 32488
rect 64390 32528 64514 32570
rect 64558 32528 64682 32570
rect 64390 32488 64392 32528
rect 64392 32488 64434 32528
rect 64434 32488 64474 32528
rect 64474 32488 64514 32528
rect 64558 32488 64598 32528
rect 64598 32488 64638 32528
rect 64638 32488 64680 32528
rect 64680 32488 64682 32528
rect 64390 32446 64514 32488
rect 64558 32446 64682 32488
rect 76390 32528 76514 32570
rect 76558 32528 76682 32570
rect 76390 32488 76392 32528
rect 76392 32488 76434 32528
rect 76434 32488 76474 32528
rect 76474 32488 76514 32528
rect 76558 32488 76598 32528
rect 76598 32488 76638 32528
rect 76638 32488 76680 32528
rect 76680 32488 76682 32528
rect 76390 32446 76514 32488
rect 76558 32446 76682 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 15150 31772 15274 31814
rect 15318 31772 15442 31814
rect 15150 31732 15152 31772
rect 15152 31732 15194 31772
rect 15194 31732 15234 31772
rect 15234 31732 15274 31772
rect 15318 31732 15358 31772
rect 15358 31732 15398 31772
rect 15398 31732 15440 31772
rect 15440 31732 15442 31772
rect 15150 31690 15274 31732
rect 15318 31690 15442 31732
rect 27150 31772 27274 31814
rect 27318 31772 27442 31814
rect 27150 31732 27152 31772
rect 27152 31732 27194 31772
rect 27194 31732 27234 31772
rect 27234 31732 27274 31772
rect 27318 31732 27358 31772
rect 27358 31732 27398 31772
rect 27398 31732 27440 31772
rect 27440 31732 27442 31772
rect 27150 31690 27274 31732
rect 27318 31690 27442 31732
rect 39150 31772 39274 31814
rect 39318 31772 39442 31814
rect 39150 31732 39152 31772
rect 39152 31732 39194 31772
rect 39194 31732 39234 31772
rect 39234 31732 39274 31772
rect 39318 31732 39358 31772
rect 39358 31732 39398 31772
rect 39398 31732 39440 31772
rect 39440 31732 39442 31772
rect 39150 31690 39274 31732
rect 39318 31690 39442 31732
rect 51150 31772 51274 31814
rect 51318 31772 51442 31814
rect 51150 31732 51152 31772
rect 51152 31732 51194 31772
rect 51194 31732 51234 31772
rect 51234 31732 51274 31772
rect 51318 31732 51358 31772
rect 51358 31732 51398 31772
rect 51398 31732 51440 31772
rect 51440 31732 51442 31772
rect 51150 31690 51274 31732
rect 51318 31690 51442 31732
rect 63150 31772 63274 31814
rect 63318 31772 63442 31814
rect 63150 31732 63152 31772
rect 63152 31732 63194 31772
rect 63194 31732 63234 31772
rect 63234 31732 63274 31772
rect 63318 31732 63358 31772
rect 63358 31732 63398 31772
rect 63398 31732 63440 31772
rect 63440 31732 63442 31772
rect 63150 31690 63274 31732
rect 63318 31690 63442 31732
rect 75150 31772 75274 31814
rect 75318 31772 75442 31814
rect 75150 31732 75152 31772
rect 75152 31732 75194 31772
rect 75194 31732 75234 31772
rect 75234 31732 75274 31772
rect 75318 31732 75358 31772
rect 75358 31732 75398 31772
rect 75398 31732 75440 31772
rect 75440 31732 75442 31772
rect 75150 31690 75274 31732
rect 75318 31690 75442 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 16390 31016 16514 31058
rect 16558 31016 16682 31058
rect 16390 30976 16392 31016
rect 16392 30976 16434 31016
rect 16434 30976 16474 31016
rect 16474 30976 16514 31016
rect 16558 30976 16598 31016
rect 16598 30976 16638 31016
rect 16638 30976 16680 31016
rect 16680 30976 16682 31016
rect 16390 30934 16514 30976
rect 16558 30934 16682 30976
rect 28390 31016 28514 31058
rect 28558 31016 28682 31058
rect 28390 30976 28392 31016
rect 28392 30976 28434 31016
rect 28434 30976 28474 31016
rect 28474 30976 28514 31016
rect 28558 30976 28598 31016
rect 28598 30976 28638 31016
rect 28638 30976 28680 31016
rect 28680 30976 28682 31016
rect 28390 30934 28514 30976
rect 28558 30934 28682 30976
rect 40390 31016 40514 31058
rect 40558 31016 40682 31058
rect 40390 30976 40392 31016
rect 40392 30976 40434 31016
rect 40434 30976 40474 31016
rect 40474 30976 40514 31016
rect 40558 30976 40598 31016
rect 40598 30976 40638 31016
rect 40638 30976 40680 31016
rect 40680 30976 40682 31016
rect 40390 30934 40514 30976
rect 40558 30934 40682 30976
rect 52390 31016 52514 31058
rect 52558 31016 52682 31058
rect 52390 30976 52392 31016
rect 52392 30976 52434 31016
rect 52434 30976 52474 31016
rect 52474 30976 52514 31016
rect 52558 30976 52598 31016
rect 52598 30976 52638 31016
rect 52638 30976 52680 31016
rect 52680 30976 52682 31016
rect 52390 30934 52514 30976
rect 52558 30934 52682 30976
rect 64390 31016 64514 31058
rect 64558 31016 64682 31058
rect 64390 30976 64392 31016
rect 64392 30976 64434 31016
rect 64434 30976 64474 31016
rect 64474 30976 64514 31016
rect 64558 30976 64598 31016
rect 64598 30976 64638 31016
rect 64638 30976 64680 31016
rect 64680 30976 64682 31016
rect 64390 30934 64514 30976
rect 64558 30934 64682 30976
rect 76390 31016 76514 31058
rect 76558 31016 76682 31058
rect 76390 30976 76392 31016
rect 76392 30976 76434 31016
rect 76434 30976 76474 31016
rect 76474 30976 76514 31016
rect 76558 30976 76598 31016
rect 76598 30976 76638 31016
rect 76638 30976 76680 31016
rect 76680 30976 76682 31016
rect 76390 30934 76514 30976
rect 76558 30934 76682 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 15150 30260 15274 30302
rect 15318 30260 15442 30302
rect 15150 30220 15152 30260
rect 15152 30220 15194 30260
rect 15194 30220 15234 30260
rect 15234 30220 15274 30260
rect 15318 30220 15358 30260
rect 15358 30220 15398 30260
rect 15398 30220 15440 30260
rect 15440 30220 15442 30260
rect 15150 30178 15274 30220
rect 15318 30178 15442 30220
rect 27150 30260 27274 30302
rect 27318 30260 27442 30302
rect 27150 30220 27152 30260
rect 27152 30220 27194 30260
rect 27194 30220 27234 30260
rect 27234 30220 27274 30260
rect 27318 30220 27358 30260
rect 27358 30220 27398 30260
rect 27398 30220 27440 30260
rect 27440 30220 27442 30260
rect 27150 30178 27274 30220
rect 27318 30178 27442 30220
rect 39150 30260 39274 30302
rect 39318 30260 39442 30302
rect 39150 30220 39152 30260
rect 39152 30220 39194 30260
rect 39194 30220 39234 30260
rect 39234 30220 39274 30260
rect 39318 30220 39358 30260
rect 39358 30220 39398 30260
rect 39398 30220 39440 30260
rect 39440 30220 39442 30260
rect 39150 30178 39274 30220
rect 39318 30178 39442 30220
rect 51150 30260 51274 30302
rect 51318 30260 51442 30302
rect 51150 30220 51152 30260
rect 51152 30220 51194 30260
rect 51194 30220 51234 30260
rect 51234 30220 51274 30260
rect 51318 30220 51358 30260
rect 51358 30220 51398 30260
rect 51398 30220 51440 30260
rect 51440 30220 51442 30260
rect 51150 30178 51274 30220
rect 51318 30178 51442 30220
rect 63150 30260 63274 30302
rect 63318 30260 63442 30302
rect 63150 30220 63152 30260
rect 63152 30220 63194 30260
rect 63194 30220 63234 30260
rect 63234 30220 63274 30260
rect 63318 30220 63358 30260
rect 63358 30220 63398 30260
rect 63398 30220 63440 30260
rect 63440 30220 63442 30260
rect 63150 30178 63274 30220
rect 63318 30178 63442 30220
rect 75150 30260 75274 30302
rect 75318 30260 75442 30302
rect 75150 30220 75152 30260
rect 75152 30220 75194 30260
rect 75194 30220 75234 30260
rect 75234 30220 75274 30260
rect 75318 30220 75358 30260
rect 75358 30220 75398 30260
rect 75398 30220 75440 30260
rect 75440 30220 75442 30260
rect 75150 30178 75274 30220
rect 75318 30178 75442 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 16390 29504 16514 29546
rect 16558 29504 16682 29546
rect 16390 29464 16392 29504
rect 16392 29464 16434 29504
rect 16434 29464 16474 29504
rect 16474 29464 16514 29504
rect 16558 29464 16598 29504
rect 16598 29464 16638 29504
rect 16638 29464 16680 29504
rect 16680 29464 16682 29504
rect 16390 29422 16514 29464
rect 16558 29422 16682 29464
rect 28390 29504 28514 29546
rect 28558 29504 28682 29546
rect 28390 29464 28392 29504
rect 28392 29464 28434 29504
rect 28434 29464 28474 29504
rect 28474 29464 28514 29504
rect 28558 29464 28598 29504
rect 28598 29464 28638 29504
rect 28638 29464 28680 29504
rect 28680 29464 28682 29504
rect 28390 29422 28514 29464
rect 28558 29422 28682 29464
rect 40390 29504 40514 29546
rect 40558 29504 40682 29546
rect 40390 29464 40392 29504
rect 40392 29464 40434 29504
rect 40434 29464 40474 29504
rect 40474 29464 40514 29504
rect 40558 29464 40598 29504
rect 40598 29464 40638 29504
rect 40638 29464 40680 29504
rect 40680 29464 40682 29504
rect 40390 29422 40514 29464
rect 40558 29422 40682 29464
rect 52390 29504 52514 29546
rect 52558 29504 52682 29546
rect 52390 29464 52392 29504
rect 52392 29464 52434 29504
rect 52434 29464 52474 29504
rect 52474 29464 52514 29504
rect 52558 29464 52598 29504
rect 52598 29464 52638 29504
rect 52638 29464 52680 29504
rect 52680 29464 52682 29504
rect 52390 29422 52514 29464
rect 52558 29422 52682 29464
rect 64390 29504 64514 29546
rect 64558 29504 64682 29546
rect 64390 29464 64392 29504
rect 64392 29464 64434 29504
rect 64434 29464 64474 29504
rect 64474 29464 64514 29504
rect 64558 29464 64598 29504
rect 64598 29464 64638 29504
rect 64638 29464 64680 29504
rect 64680 29464 64682 29504
rect 64390 29422 64514 29464
rect 64558 29422 64682 29464
rect 76390 29504 76514 29546
rect 76558 29504 76682 29546
rect 76390 29464 76392 29504
rect 76392 29464 76434 29504
rect 76434 29464 76474 29504
rect 76474 29464 76514 29504
rect 76558 29464 76598 29504
rect 76598 29464 76638 29504
rect 76638 29464 76680 29504
rect 76680 29464 76682 29504
rect 76390 29422 76514 29464
rect 76558 29422 76682 29464
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 15150 28748 15274 28790
rect 15318 28748 15442 28790
rect 15150 28708 15152 28748
rect 15152 28708 15194 28748
rect 15194 28708 15234 28748
rect 15234 28708 15274 28748
rect 15318 28708 15358 28748
rect 15358 28708 15398 28748
rect 15398 28708 15440 28748
rect 15440 28708 15442 28748
rect 15150 28666 15274 28708
rect 15318 28666 15442 28708
rect 27150 28748 27274 28790
rect 27318 28748 27442 28790
rect 27150 28708 27152 28748
rect 27152 28708 27194 28748
rect 27194 28708 27234 28748
rect 27234 28708 27274 28748
rect 27318 28708 27358 28748
rect 27358 28708 27398 28748
rect 27398 28708 27440 28748
rect 27440 28708 27442 28748
rect 27150 28666 27274 28708
rect 27318 28666 27442 28708
rect 39150 28748 39274 28790
rect 39318 28748 39442 28790
rect 39150 28708 39152 28748
rect 39152 28708 39194 28748
rect 39194 28708 39234 28748
rect 39234 28708 39274 28748
rect 39318 28708 39358 28748
rect 39358 28708 39398 28748
rect 39398 28708 39440 28748
rect 39440 28708 39442 28748
rect 39150 28666 39274 28708
rect 39318 28666 39442 28708
rect 51150 28748 51274 28790
rect 51318 28748 51442 28790
rect 51150 28708 51152 28748
rect 51152 28708 51194 28748
rect 51194 28708 51234 28748
rect 51234 28708 51274 28748
rect 51318 28708 51358 28748
rect 51358 28708 51398 28748
rect 51398 28708 51440 28748
rect 51440 28708 51442 28748
rect 51150 28666 51274 28708
rect 51318 28666 51442 28708
rect 63150 28748 63274 28790
rect 63318 28748 63442 28790
rect 63150 28708 63152 28748
rect 63152 28708 63194 28748
rect 63194 28708 63234 28748
rect 63234 28708 63274 28748
rect 63318 28708 63358 28748
rect 63358 28708 63398 28748
rect 63398 28708 63440 28748
rect 63440 28708 63442 28748
rect 63150 28666 63274 28708
rect 63318 28666 63442 28708
rect 75150 28748 75274 28790
rect 75318 28748 75442 28790
rect 75150 28708 75152 28748
rect 75152 28708 75194 28748
rect 75194 28708 75234 28748
rect 75234 28708 75274 28748
rect 75318 28708 75358 28748
rect 75358 28708 75398 28748
rect 75398 28708 75440 28748
rect 75440 28708 75442 28748
rect 75150 28666 75274 28708
rect 75318 28666 75442 28708
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 16390 27992 16514 28034
rect 16558 27992 16682 28034
rect 16390 27952 16392 27992
rect 16392 27952 16434 27992
rect 16434 27952 16474 27992
rect 16474 27952 16514 27992
rect 16558 27952 16598 27992
rect 16598 27952 16638 27992
rect 16638 27952 16680 27992
rect 16680 27952 16682 27992
rect 16390 27910 16514 27952
rect 16558 27910 16682 27952
rect 28390 27992 28514 28034
rect 28558 27992 28682 28034
rect 28390 27952 28392 27992
rect 28392 27952 28434 27992
rect 28434 27952 28474 27992
rect 28474 27952 28514 27992
rect 28558 27952 28598 27992
rect 28598 27952 28638 27992
rect 28638 27952 28680 27992
rect 28680 27952 28682 27992
rect 28390 27910 28514 27952
rect 28558 27910 28682 27952
rect 40390 27992 40514 28034
rect 40558 27992 40682 28034
rect 40390 27952 40392 27992
rect 40392 27952 40434 27992
rect 40434 27952 40474 27992
rect 40474 27952 40514 27992
rect 40558 27952 40598 27992
rect 40598 27952 40638 27992
rect 40638 27952 40680 27992
rect 40680 27952 40682 27992
rect 40390 27910 40514 27952
rect 40558 27910 40682 27952
rect 52390 27992 52514 28034
rect 52558 27992 52682 28034
rect 52390 27952 52392 27992
rect 52392 27952 52434 27992
rect 52434 27952 52474 27992
rect 52474 27952 52514 27992
rect 52558 27952 52598 27992
rect 52598 27952 52638 27992
rect 52638 27952 52680 27992
rect 52680 27952 52682 27992
rect 52390 27910 52514 27952
rect 52558 27910 52682 27952
rect 64390 27992 64514 28034
rect 64558 27992 64682 28034
rect 64390 27952 64392 27992
rect 64392 27952 64434 27992
rect 64434 27952 64474 27992
rect 64474 27952 64514 27992
rect 64558 27952 64598 27992
rect 64598 27952 64638 27992
rect 64638 27952 64680 27992
rect 64680 27952 64682 27992
rect 64390 27910 64514 27952
rect 64558 27910 64682 27952
rect 76390 27992 76514 28034
rect 76558 27992 76682 28034
rect 76390 27952 76392 27992
rect 76392 27952 76434 27992
rect 76434 27952 76474 27992
rect 76474 27952 76514 27992
rect 76558 27952 76598 27992
rect 76598 27952 76638 27992
rect 76638 27952 76680 27992
rect 76680 27952 76682 27992
rect 76390 27910 76514 27952
rect 76558 27910 76682 27952
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 15150 27236 15274 27278
rect 15318 27236 15442 27278
rect 15150 27196 15152 27236
rect 15152 27196 15194 27236
rect 15194 27196 15234 27236
rect 15234 27196 15274 27236
rect 15318 27196 15358 27236
rect 15358 27196 15398 27236
rect 15398 27196 15440 27236
rect 15440 27196 15442 27236
rect 15150 27154 15274 27196
rect 15318 27154 15442 27196
rect 27150 27236 27274 27278
rect 27318 27236 27442 27278
rect 27150 27196 27152 27236
rect 27152 27196 27194 27236
rect 27194 27196 27234 27236
rect 27234 27196 27274 27236
rect 27318 27196 27358 27236
rect 27358 27196 27398 27236
rect 27398 27196 27440 27236
rect 27440 27196 27442 27236
rect 27150 27154 27274 27196
rect 27318 27154 27442 27196
rect 39150 27236 39274 27278
rect 39318 27236 39442 27278
rect 39150 27196 39152 27236
rect 39152 27196 39194 27236
rect 39194 27196 39234 27236
rect 39234 27196 39274 27236
rect 39318 27196 39358 27236
rect 39358 27196 39398 27236
rect 39398 27196 39440 27236
rect 39440 27196 39442 27236
rect 39150 27154 39274 27196
rect 39318 27154 39442 27196
rect 51150 27236 51274 27278
rect 51318 27236 51442 27278
rect 51150 27196 51152 27236
rect 51152 27196 51194 27236
rect 51194 27196 51234 27236
rect 51234 27196 51274 27236
rect 51318 27196 51358 27236
rect 51358 27196 51398 27236
rect 51398 27196 51440 27236
rect 51440 27196 51442 27236
rect 51150 27154 51274 27196
rect 51318 27154 51442 27196
rect 63150 27236 63274 27278
rect 63318 27236 63442 27278
rect 63150 27196 63152 27236
rect 63152 27196 63194 27236
rect 63194 27196 63234 27236
rect 63234 27196 63274 27236
rect 63318 27196 63358 27236
rect 63358 27196 63398 27236
rect 63398 27196 63440 27236
rect 63440 27196 63442 27236
rect 63150 27154 63274 27196
rect 63318 27154 63442 27196
rect 75150 27236 75274 27278
rect 75318 27236 75442 27278
rect 75150 27196 75152 27236
rect 75152 27196 75194 27236
rect 75194 27196 75234 27236
rect 75234 27196 75274 27236
rect 75318 27196 75358 27236
rect 75358 27196 75398 27236
rect 75398 27196 75440 27236
rect 75440 27196 75442 27236
rect 75150 27154 75274 27196
rect 75318 27154 75442 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 16390 26480 16514 26522
rect 16558 26480 16682 26522
rect 16390 26440 16392 26480
rect 16392 26440 16434 26480
rect 16434 26440 16474 26480
rect 16474 26440 16514 26480
rect 16558 26440 16598 26480
rect 16598 26440 16638 26480
rect 16638 26440 16680 26480
rect 16680 26440 16682 26480
rect 16390 26398 16514 26440
rect 16558 26398 16682 26440
rect 28390 26480 28514 26522
rect 28558 26480 28682 26522
rect 28390 26440 28392 26480
rect 28392 26440 28434 26480
rect 28434 26440 28474 26480
rect 28474 26440 28514 26480
rect 28558 26440 28598 26480
rect 28598 26440 28638 26480
rect 28638 26440 28680 26480
rect 28680 26440 28682 26480
rect 28390 26398 28514 26440
rect 28558 26398 28682 26440
rect 40390 26480 40514 26522
rect 40558 26480 40682 26522
rect 40390 26440 40392 26480
rect 40392 26440 40434 26480
rect 40434 26440 40474 26480
rect 40474 26440 40514 26480
rect 40558 26440 40598 26480
rect 40598 26440 40638 26480
rect 40638 26440 40680 26480
rect 40680 26440 40682 26480
rect 40390 26398 40514 26440
rect 40558 26398 40682 26440
rect 52390 26480 52514 26522
rect 52558 26480 52682 26522
rect 64390 26480 64514 26522
rect 64558 26480 64682 26522
rect 52390 26440 52392 26480
rect 52392 26440 52434 26480
rect 52434 26440 52474 26480
rect 52474 26440 52514 26480
rect 52558 26440 52598 26480
rect 52598 26440 52638 26480
rect 52638 26440 52680 26480
rect 52680 26440 52682 26480
rect 64390 26440 64392 26480
rect 64392 26440 64434 26480
rect 64434 26440 64474 26480
rect 64474 26440 64514 26480
rect 64558 26440 64598 26480
rect 64598 26440 64638 26480
rect 64638 26440 64680 26480
rect 64680 26440 64682 26480
rect 52390 26398 52514 26440
rect 52558 26398 52682 26440
rect 64390 26398 64514 26440
rect 64558 26398 64682 26440
rect 76390 26480 76514 26522
rect 76558 26480 76682 26522
rect 76390 26440 76392 26480
rect 76392 26440 76434 26480
rect 76434 26440 76474 26480
rect 76474 26440 76514 26480
rect 76558 26440 76598 26480
rect 76598 26440 76638 26480
rect 76638 26440 76680 26480
rect 76680 26440 76682 26480
rect 76390 26398 76514 26440
rect 76558 26398 76682 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 15150 25724 15274 25766
rect 15318 25724 15442 25766
rect 15150 25684 15152 25724
rect 15152 25684 15194 25724
rect 15194 25684 15234 25724
rect 15234 25684 15274 25724
rect 15318 25684 15358 25724
rect 15358 25684 15398 25724
rect 15398 25684 15440 25724
rect 15440 25684 15442 25724
rect 15150 25642 15274 25684
rect 15318 25642 15442 25684
rect 27150 25724 27274 25766
rect 27318 25724 27442 25766
rect 27150 25684 27152 25724
rect 27152 25684 27194 25724
rect 27194 25684 27234 25724
rect 27234 25684 27274 25724
rect 27318 25684 27358 25724
rect 27358 25684 27398 25724
rect 27398 25684 27440 25724
rect 27440 25684 27442 25724
rect 27150 25642 27274 25684
rect 27318 25642 27442 25684
rect 39150 25724 39274 25766
rect 39318 25724 39442 25766
rect 39150 25684 39152 25724
rect 39152 25684 39194 25724
rect 39194 25684 39234 25724
rect 39234 25684 39274 25724
rect 39318 25684 39358 25724
rect 39358 25684 39398 25724
rect 39398 25684 39440 25724
rect 39440 25684 39442 25724
rect 39150 25642 39274 25684
rect 39318 25642 39442 25684
rect 51150 25724 51274 25766
rect 51318 25724 51442 25766
rect 51150 25684 51152 25724
rect 51152 25684 51194 25724
rect 51194 25684 51234 25724
rect 51234 25684 51274 25724
rect 51318 25684 51358 25724
rect 51358 25684 51398 25724
rect 51398 25684 51440 25724
rect 51440 25684 51442 25724
rect 51150 25642 51274 25684
rect 51318 25642 51442 25684
rect 63150 25724 63274 25766
rect 63318 25724 63442 25766
rect 63150 25684 63152 25724
rect 63152 25684 63194 25724
rect 63194 25684 63234 25724
rect 63234 25684 63274 25724
rect 63318 25684 63358 25724
rect 63358 25684 63398 25724
rect 63398 25684 63440 25724
rect 63440 25684 63442 25724
rect 63150 25642 63274 25684
rect 63318 25642 63442 25684
rect 75150 25724 75274 25766
rect 75318 25724 75442 25766
rect 75150 25684 75152 25724
rect 75152 25684 75194 25724
rect 75194 25684 75234 25724
rect 75234 25684 75274 25724
rect 75318 25684 75358 25724
rect 75358 25684 75398 25724
rect 75398 25684 75440 25724
rect 75440 25684 75442 25724
rect 75150 25642 75274 25684
rect 75318 25642 75442 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 16390 24968 16514 25010
rect 16558 24968 16682 25010
rect 16390 24928 16392 24968
rect 16392 24928 16434 24968
rect 16434 24928 16474 24968
rect 16474 24928 16514 24968
rect 16558 24928 16598 24968
rect 16598 24928 16638 24968
rect 16638 24928 16680 24968
rect 16680 24928 16682 24968
rect 16390 24886 16514 24928
rect 16558 24886 16682 24928
rect 28390 24968 28514 25010
rect 28558 24968 28682 25010
rect 28390 24928 28392 24968
rect 28392 24928 28434 24968
rect 28434 24928 28474 24968
rect 28474 24928 28514 24968
rect 28558 24928 28598 24968
rect 28598 24928 28638 24968
rect 28638 24928 28680 24968
rect 28680 24928 28682 24968
rect 28390 24886 28514 24928
rect 28558 24886 28682 24928
rect 40390 24968 40514 25010
rect 40558 24968 40682 25010
rect 40390 24928 40392 24968
rect 40392 24928 40434 24968
rect 40434 24928 40474 24968
rect 40474 24928 40514 24968
rect 40558 24928 40598 24968
rect 40598 24928 40638 24968
rect 40638 24928 40680 24968
rect 40680 24928 40682 24968
rect 40390 24886 40514 24928
rect 40558 24886 40682 24928
rect 52390 24968 52514 25010
rect 52558 24968 52682 25010
rect 52390 24928 52392 24968
rect 52392 24928 52434 24968
rect 52434 24928 52474 24968
rect 52474 24928 52514 24968
rect 52558 24928 52598 24968
rect 52598 24928 52638 24968
rect 52638 24928 52680 24968
rect 52680 24928 52682 24968
rect 52390 24886 52514 24928
rect 52558 24886 52682 24928
rect 64390 24968 64514 25010
rect 64558 24968 64682 25010
rect 64390 24928 64392 24968
rect 64392 24928 64434 24968
rect 64434 24928 64474 24968
rect 64474 24928 64514 24968
rect 64558 24928 64598 24968
rect 64598 24928 64638 24968
rect 64638 24928 64680 24968
rect 64680 24928 64682 24968
rect 64390 24886 64514 24928
rect 64558 24886 64682 24928
rect 76390 24968 76514 25010
rect 76558 24968 76682 25010
rect 76390 24928 76392 24968
rect 76392 24928 76434 24968
rect 76434 24928 76474 24968
rect 76474 24928 76514 24968
rect 76558 24928 76598 24968
rect 76598 24928 76638 24968
rect 76638 24928 76680 24968
rect 76680 24928 76682 24968
rect 76390 24886 76514 24928
rect 76558 24886 76682 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 15150 24212 15274 24254
rect 15318 24212 15442 24254
rect 15150 24172 15152 24212
rect 15152 24172 15194 24212
rect 15194 24172 15234 24212
rect 15234 24172 15274 24212
rect 15318 24172 15358 24212
rect 15358 24172 15398 24212
rect 15398 24172 15440 24212
rect 15440 24172 15442 24212
rect 15150 24130 15274 24172
rect 15318 24130 15442 24172
rect 27150 24212 27274 24254
rect 27318 24212 27442 24254
rect 27150 24172 27152 24212
rect 27152 24172 27194 24212
rect 27194 24172 27234 24212
rect 27234 24172 27274 24212
rect 27318 24172 27358 24212
rect 27358 24172 27398 24212
rect 27398 24172 27440 24212
rect 27440 24172 27442 24212
rect 27150 24130 27274 24172
rect 27318 24130 27442 24172
rect 39150 24212 39274 24254
rect 39318 24212 39442 24254
rect 39150 24172 39152 24212
rect 39152 24172 39194 24212
rect 39194 24172 39234 24212
rect 39234 24172 39274 24212
rect 39318 24172 39358 24212
rect 39358 24172 39398 24212
rect 39398 24172 39440 24212
rect 39440 24172 39442 24212
rect 39150 24130 39274 24172
rect 39318 24130 39442 24172
rect 78698 23710 78822 23834
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 16390 23456 16514 23498
rect 16558 23456 16682 23498
rect 16390 23416 16392 23456
rect 16392 23416 16434 23456
rect 16434 23416 16474 23456
rect 16474 23416 16514 23456
rect 16558 23416 16598 23456
rect 16598 23416 16638 23456
rect 16638 23416 16680 23456
rect 16680 23416 16682 23456
rect 16390 23374 16514 23416
rect 16558 23374 16682 23416
rect 28390 23456 28514 23498
rect 28558 23456 28682 23498
rect 28390 23416 28392 23456
rect 28392 23416 28434 23456
rect 28434 23416 28474 23456
rect 28474 23416 28514 23456
rect 28558 23416 28598 23456
rect 28598 23416 28638 23456
rect 28638 23416 28680 23456
rect 28680 23416 28682 23456
rect 28390 23374 28514 23416
rect 28558 23374 28682 23416
rect 40390 23456 40514 23498
rect 40558 23456 40682 23498
rect 40390 23416 40392 23456
rect 40392 23416 40434 23456
rect 40434 23416 40474 23456
rect 40474 23416 40514 23456
rect 40558 23416 40598 23456
rect 40598 23416 40638 23456
rect 40638 23416 40680 23456
rect 40680 23416 40682 23456
rect 40390 23374 40514 23416
rect 40558 23374 40682 23416
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 15150 22700 15274 22742
rect 15318 22700 15442 22742
rect 15150 22660 15152 22700
rect 15152 22660 15194 22700
rect 15194 22660 15234 22700
rect 15234 22660 15274 22700
rect 15318 22660 15358 22700
rect 15358 22660 15398 22700
rect 15398 22660 15440 22700
rect 15440 22660 15442 22700
rect 15150 22618 15274 22660
rect 15318 22618 15442 22660
rect 27150 22700 27274 22742
rect 27318 22700 27442 22742
rect 27150 22660 27152 22700
rect 27152 22660 27194 22700
rect 27194 22660 27234 22700
rect 27234 22660 27274 22700
rect 27318 22660 27358 22700
rect 27358 22660 27398 22700
rect 27398 22660 27440 22700
rect 27440 22660 27442 22700
rect 27150 22618 27274 22660
rect 27318 22618 27442 22660
rect 39150 22700 39274 22742
rect 39318 22700 39442 22742
rect 39150 22660 39152 22700
rect 39152 22660 39194 22700
rect 39194 22660 39234 22700
rect 39234 22660 39274 22700
rect 39318 22660 39358 22700
rect 39358 22660 39398 22700
rect 39398 22660 39440 22700
rect 39440 22660 39442 22700
rect 39150 22618 39274 22660
rect 39318 22618 39442 22660
rect 64390 22417 64514 22541
rect 64558 22417 64682 22541
rect 64390 22249 64514 22373
rect 64558 22249 64682 22373
rect 64390 22081 64514 22205
rect 64558 22081 64682 22205
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 16390 21944 16514 21986
rect 16558 21944 16682 21986
rect 16390 21904 16392 21944
rect 16392 21904 16434 21944
rect 16434 21904 16474 21944
rect 16474 21904 16514 21944
rect 16558 21904 16598 21944
rect 16598 21904 16638 21944
rect 16638 21904 16680 21944
rect 16680 21904 16682 21944
rect 16390 21862 16514 21904
rect 16558 21862 16682 21904
rect 28390 21944 28514 21986
rect 28558 21944 28682 21986
rect 28390 21904 28392 21944
rect 28392 21904 28434 21944
rect 28434 21904 28474 21944
rect 28474 21904 28514 21944
rect 28558 21904 28598 21944
rect 28598 21904 28638 21944
rect 28638 21904 28680 21944
rect 28680 21904 28682 21944
rect 28390 21862 28514 21904
rect 28558 21862 28682 21904
rect 40390 21944 40514 21986
rect 40558 21944 40682 21986
rect 40390 21904 40392 21944
rect 40392 21904 40434 21944
rect 40434 21904 40474 21944
rect 40474 21904 40514 21944
rect 40558 21904 40598 21944
rect 40598 21904 40638 21944
rect 40638 21904 40680 21944
rect 40680 21904 40682 21944
rect 40390 21862 40514 21904
rect 40558 21862 40682 21904
rect 64390 21913 64514 22037
rect 64558 21913 64682 22037
rect 64390 21745 64514 21869
rect 64558 21745 64682 21869
rect 64390 21577 64514 21701
rect 64558 21577 64682 21701
rect 64390 21409 64514 21533
rect 64558 21409 64682 21533
rect 64390 21241 64514 21365
rect 64558 21241 64682 21365
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 15150 21188 15274 21230
rect 15318 21188 15442 21230
rect 15150 21148 15152 21188
rect 15152 21148 15194 21188
rect 15194 21148 15234 21188
rect 15234 21148 15274 21188
rect 15318 21148 15358 21188
rect 15358 21148 15398 21188
rect 15398 21148 15440 21188
rect 15440 21148 15442 21188
rect 15150 21106 15274 21148
rect 15318 21106 15442 21148
rect 27150 21188 27274 21230
rect 27318 21188 27442 21230
rect 27150 21148 27152 21188
rect 27152 21148 27194 21188
rect 27194 21148 27234 21188
rect 27234 21148 27274 21188
rect 27318 21148 27358 21188
rect 27358 21148 27398 21188
rect 27398 21148 27440 21188
rect 27440 21148 27442 21188
rect 27150 21106 27274 21148
rect 27318 21106 27442 21148
rect 39150 21188 39274 21230
rect 39318 21188 39442 21230
rect 39150 21148 39152 21188
rect 39152 21148 39194 21188
rect 39194 21148 39234 21188
rect 39234 21148 39274 21188
rect 39318 21148 39358 21188
rect 39358 21148 39398 21188
rect 39398 21148 39440 21188
rect 39440 21148 39442 21188
rect 39150 21106 39274 21148
rect 39318 21106 39442 21148
rect 64390 21073 64514 21197
rect 64558 21073 64682 21197
rect 64390 20905 64514 21029
rect 64558 20905 64682 21029
rect 64390 20737 64514 20861
rect 64558 20737 64682 20861
rect 64390 20569 64514 20693
rect 64558 20569 64682 20693
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 16390 20432 16514 20474
rect 16558 20432 16682 20474
rect 16390 20392 16392 20432
rect 16392 20392 16434 20432
rect 16434 20392 16474 20432
rect 16474 20392 16514 20432
rect 16558 20392 16598 20432
rect 16598 20392 16638 20432
rect 16638 20392 16680 20432
rect 16680 20392 16682 20432
rect 16390 20350 16514 20392
rect 16558 20350 16682 20392
rect 28390 20432 28514 20474
rect 28558 20432 28682 20474
rect 28390 20392 28392 20432
rect 28392 20392 28434 20432
rect 28434 20392 28474 20432
rect 28474 20392 28514 20432
rect 28558 20392 28598 20432
rect 28598 20392 28638 20432
rect 28638 20392 28680 20432
rect 28680 20392 28682 20432
rect 28390 20350 28514 20392
rect 28558 20350 28682 20392
rect 40390 20432 40514 20474
rect 40558 20432 40682 20474
rect 40390 20392 40392 20432
rect 40392 20392 40434 20432
rect 40434 20392 40474 20432
rect 40474 20392 40514 20432
rect 40558 20392 40598 20432
rect 40598 20392 40638 20432
rect 40638 20392 40680 20432
rect 40680 20392 40682 20432
rect 40390 20350 40514 20392
rect 40558 20350 40682 20392
rect 64390 20401 64514 20525
rect 64558 20401 64682 20525
rect 76390 22417 76514 22541
rect 76558 22417 76682 22541
rect 76390 22249 76514 22373
rect 76558 22249 76682 22373
rect 76390 22081 76514 22205
rect 76558 22081 76682 22205
rect 76390 21913 76514 22037
rect 76558 21913 76682 22037
rect 76390 21745 76514 21869
rect 76558 21745 76682 21869
rect 76390 21577 76514 21701
rect 76558 21577 76682 21701
rect 76390 21409 76514 21533
rect 76558 21409 76682 21533
rect 76390 21241 76514 21365
rect 76558 21241 76682 21365
rect 76390 21073 76514 21197
rect 76558 21073 76682 21197
rect 76390 20905 76514 21029
rect 76558 20905 76682 21029
rect 76390 20737 76514 20861
rect 76558 20737 76682 20861
rect 76390 20569 76514 20693
rect 76558 20569 76682 20693
rect 76390 20401 76514 20525
rect 76558 20401 76682 20525
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 15150 19676 15274 19718
rect 15318 19676 15442 19718
rect 15150 19636 15152 19676
rect 15152 19636 15194 19676
rect 15194 19636 15234 19676
rect 15234 19636 15274 19676
rect 15318 19636 15358 19676
rect 15358 19636 15398 19676
rect 15398 19636 15440 19676
rect 15440 19636 15442 19676
rect 15150 19594 15274 19636
rect 15318 19594 15442 19636
rect 27150 19676 27274 19718
rect 27318 19676 27442 19718
rect 27150 19636 27152 19676
rect 27152 19636 27194 19676
rect 27194 19636 27234 19676
rect 27234 19636 27274 19676
rect 27318 19636 27358 19676
rect 27358 19636 27398 19676
rect 27398 19636 27440 19676
rect 27440 19636 27442 19676
rect 27150 19594 27274 19636
rect 27318 19594 27442 19636
rect 39150 19676 39274 19718
rect 39318 19676 39442 19718
rect 39150 19636 39152 19676
rect 39152 19636 39194 19676
rect 39194 19636 39234 19676
rect 39234 19636 39274 19676
rect 39318 19636 39358 19676
rect 39358 19636 39398 19676
rect 39398 19636 39440 19676
rect 39440 19636 39442 19676
rect 39150 19594 39274 19636
rect 39318 19594 39442 19636
rect 63150 19541 63274 19665
rect 63318 19541 63442 19665
rect 63150 19373 63274 19497
rect 63318 19373 63442 19497
rect 63150 19205 63274 19329
rect 63318 19205 63442 19329
rect 63150 19037 63274 19161
rect 63318 19037 63442 19161
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 16390 18920 16514 18962
rect 16558 18920 16682 18962
rect 16390 18880 16392 18920
rect 16392 18880 16434 18920
rect 16434 18880 16474 18920
rect 16474 18880 16514 18920
rect 16558 18880 16598 18920
rect 16598 18880 16638 18920
rect 16638 18880 16680 18920
rect 16680 18880 16682 18920
rect 16390 18838 16514 18880
rect 16558 18838 16682 18880
rect 28390 18920 28514 18962
rect 28558 18920 28682 18962
rect 28390 18880 28392 18920
rect 28392 18880 28434 18920
rect 28434 18880 28474 18920
rect 28474 18880 28514 18920
rect 28558 18880 28598 18920
rect 28598 18880 28638 18920
rect 28638 18880 28680 18920
rect 28680 18880 28682 18920
rect 28390 18838 28514 18880
rect 28558 18838 28682 18880
rect 40390 18920 40514 18962
rect 40558 18920 40682 18962
rect 40390 18880 40392 18920
rect 40392 18880 40434 18920
rect 40434 18880 40474 18920
rect 40474 18880 40514 18920
rect 40558 18880 40598 18920
rect 40598 18880 40638 18920
rect 40638 18880 40680 18920
rect 40680 18880 40682 18920
rect 40390 18838 40514 18880
rect 40558 18838 40682 18880
rect 63150 18869 63274 18993
rect 63318 18869 63442 18993
rect 63150 18701 63274 18825
rect 63318 18701 63442 18825
rect 63150 18533 63274 18657
rect 63318 18533 63442 18657
rect 63150 18365 63274 18489
rect 63318 18365 63442 18489
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 15150 18164 15274 18206
rect 15318 18164 15442 18206
rect 15150 18124 15152 18164
rect 15152 18124 15194 18164
rect 15194 18124 15234 18164
rect 15234 18124 15274 18164
rect 15318 18124 15358 18164
rect 15358 18124 15398 18164
rect 15398 18124 15440 18164
rect 15440 18124 15442 18164
rect 15150 18082 15274 18124
rect 15318 18082 15442 18124
rect 27150 18164 27274 18206
rect 27318 18164 27442 18206
rect 27150 18124 27152 18164
rect 27152 18124 27194 18164
rect 27194 18124 27234 18164
rect 27234 18124 27274 18164
rect 27318 18124 27358 18164
rect 27358 18124 27398 18164
rect 27398 18124 27440 18164
rect 27440 18124 27442 18164
rect 27150 18082 27274 18124
rect 27318 18082 27442 18124
rect 39150 18164 39274 18206
rect 39318 18164 39442 18206
rect 39150 18124 39152 18164
rect 39152 18124 39194 18164
rect 39194 18124 39234 18164
rect 39234 18124 39274 18164
rect 39318 18124 39358 18164
rect 39358 18124 39398 18164
rect 39398 18124 39440 18164
rect 39440 18124 39442 18164
rect 39150 18082 39274 18124
rect 39318 18082 39442 18124
rect 63150 18197 63274 18321
rect 63318 18197 63442 18321
rect 63150 18029 63274 18153
rect 63318 18029 63442 18153
rect 63150 17861 63274 17985
rect 63318 17861 63442 17985
rect 63150 17693 63274 17817
rect 63318 17693 63442 17817
rect 63150 17525 63274 17649
rect 63318 17525 63442 17649
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 16390 17408 16514 17450
rect 16558 17408 16682 17450
rect 16390 17368 16392 17408
rect 16392 17368 16434 17408
rect 16434 17368 16474 17408
rect 16474 17368 16514 17408
rect 16558 17368 16598 17408
rect 16598 17368 16638 17408
rect 16638 17368 16680 17408
rect 16680 17368 16682 17408
rect 16390 17326 16514 17368
rect 16558 17326 16682 17368
rect 28390 17408 28514 17450
rect 28558 17408 28682 17450
rect 28390 17368 28392 17408
rect 28392 17368 28434 17408
rect 28434 17368 28474 17408
rect 28474 17368 28514 17408
rect 28558 17368 28598 17408
rect 28598 17368 28638 17408
rect 28638 17368 28680 17408
rect 28680 17368 28682 17408
rect 28390 17326 28514 17368
rect 28558 17326 28682 17368
rect 40390 17408 40514 17450
rect 40558 17408 40682 17450
rect 75150 19541 75274 19665
rect 75318 19541 75442 19665
rect 75150 19373 75274 19497
rect 75318 19373 75442 19497
rect 75150 19205 75274 19329
rect 75318 19205 75442 19329
rect 75150 19037 75274 19161
rect 75318 19037 75442 19161
rect 75150 18869 75274 18993
rect 75318 18869 75442 18993
rect 75150 18701 75274 18825
rect 75318 18701 75442 18825
rect 75150 18533 75274 18657
rect 75318 18533 75442 18657
rect 75150 18365 75274 18489
rect 75318 18365 75442 18489
rect 75150 18197 75274 18321
rect 75318 18197 75442 18321
rect 75150 18029 75274 18153
rect 75318 18029 75442 18153
rect 75150 17861 75274 17985
rect 75318 17861 75442 17985
rect 75150 17693 75274 17817
rect 75318 17693 75442 17817
rect 75150 17525 75274 17649
rect 75318 17525 75442 17649
rect 40390 17368 40392 17408
rect 40392 17368 40434 17408
rect 40434 17368 40474 17408
rect 40474 17368 40514 17408
rect 40558 17368 40598 17408
rect 40598 17368 40638 17408
rect 40638 17368 40680 17408
rect 40680 17368 40682 17408
rect 40390 17326 40514 17368
rect 40558 17326 40682 17368
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 15150 16652 15274 16694
rect 15318 16652 15442 16694
rect 15150 16612 15152 16652
rect 15152 16612 15194 16652
rect 15194 16612 15234 16652
rect 15234 16612 15274 16652
rect 15318 16612 15358 16652
rect 15358 16612 15398 16652
rect 15398 16612 15440 16652
rect 15440 16612 15442 16652
rect 15150 16570 15274 16612
rect 15318 16570 15442 16612
rect 27150 16652 27274 16694
rect 27318 16652 27442 16694
rect 27150 16612 27152 16652
rect 27152 16612 27194 16652
rect 27194 16612 27234 16652
rect 27234 16612 27274 16652
rect 27318 16612 27358 16652
rect 27358 16612 27398 16652
rect 27398 16612 27440 16652
rect 27440 16612 27442 16652
rect 27150 16570 27274 16612
rect 27318 16570 27442 16612
rect 39150 16652 39274 16694
rect 39318 16652 39442 16694
rect 39150 16612 39152 16652
rect 39152 16612 39194 16652
rect 39194 16612 39234 16652
rect 39234 16612 39274 16652
rect 39318 16612 39358 16652
rect 39358 16612 39398 16652
rect 39398 16612 39440 16652
rect 39440 16612 39442 16652
rect 39150 16570 39274 16612
rect 39318 16570 39442 16612
rect 78698 16150 78822 16274
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 16390 15896 16514 15938
rect 16558 15896 16682 15938
rect 16390 15856 16392 15896
rect 16392 15856 16434 15896
rect 16434 15856 16474 15896
rect 16474 15856 16514 15896
rect 16558 15856 16598 15896
rect 16598 15856 16638 15896
rect 16638 15856 16680 15896
rect 16680 15856 16682 15896
rect 16390 15814 16514 15856
rect 16558 15814 16682 15856
rect 28390 15896 28514 15938
rect 28558 15896 28682 15938
rect 28390 15856 28392 15896
rect 28392 15856 28434 15896
rect 28434 15856 28474 15896
rect 28474 15856 28514 15896
rect 28558 15856 28598 15896
rect 28598 15856 28638 15896
rect 28638 15856 28680 15896
rect 28680 15856 28682 15896
rect 28390 15814 28514 15856
rect 28558 15814 28682 15856
rect 40390 15896 40514 15938
rect 40558 15896 40682 15938
rect 40390 15856 40392 15896
rect 40392 15856 40434 15896
rect 40434 15856 40474 15896
rect 40474 15856 40514 15896
rect 40558 15856 40598 15896
rect 40598 15856 40638 15896
rect 40638 15856 40680 15896
rect 40680 15856 40682 15896
rect 40390 15814 40514 15856
rect 40558 15814 40682 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 15150 15140 15274 15182
rect 15318 15140 15442 15182
rect 15150 15100 15152 15140
rect 15152 15100 15194 15140
rect 15194 15100 15234 15140
rect 15234 15100 15274 15140
rect 15318 15100 15358 15140
rect 15358 15100 15398 15140
rect 15398 15100 15440 15140
rect 15440 15100 15442 15140
rect 15150 15058 15274 15100
rect 15318 15058 15442 15100
rect 27150 15140 27274 15182
rect 27318 15140 27442 15182
rect 27150 15100 27152 15140
rect 27152 15100 27194 15140
rect 27194 15100 27234 15140
rect 27234 15100 27274 15140
rect 27318 15100 27358 15140
rect 27358 15100 27398 15140
rect 27398 15100 27440 15140
rect 27440 15100 27442 15140
rect 27150 15058 27274 15100
rect 27318 15058 27442 15100
rect 39150 15140 39274 15182
rect 39318 15140 39442 15182
rect 39150 15100 39152 15140
rect 39152 15100 39194 15140
rect 39194 15100 39234 15140
rect 39234 15100 39274 15140
rect 39318 15100 39358 15140
rect 39358 15100 39398 15140
rect 39398 15100 39440 15140
rect 39440 15100 39442 15140
rect 39150 15058 39274 15100
rect 39318 15058 39442 15100
rect 51150 15140 51274 15182
rect 51318 15140 51442 15182
rect 51150 15100 51152 15140
rect 51152 15100 51194 15140
rect 51194 15100 51234 15140
rect 51234 15100 51274 15140
rect 51318 15100 51358 15140
rect 51358 15100 51398 15140
rect 51398 15100 51440 15140
rect 51440 15100 51442 15140
rect 51150 15058 51274 15100
rect 51318 15058 51442 15100
rect 63150 15140 63274 15182
rect 63318 15140 63442 15182
rect 63150 15100 63152 15140
rect 63152 15100 63194 15140
rect 63194 15100 63234 15140
rect 63234 15100 63274 15140
rect 63318 15100 63358 15140
rect 63358 15100 63398 15140
rect 63398 15100 63440 15140
rect 63440 15100 63442 15140
rect 63150 15058 63274 15100
rect 63318 15058 63442 15100
rect 75150 15140 75274 15182
rect 75318 15140 75442 15182
rect 75150 15100 75152 15140
rect 75152 15100 75194 15140
rect 75194 15100 75234 15140
rect 75234 15100 75274 15140
rect 75318 15100 75358 15140
rect 75358 15100 75398 15140
rect 75398 15100 75440 15140
rect 75440 15100 75442 15140
rect 75150 15058 75274 15100
rect 75318 15058 75442 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 16390 14384 16514 14426
rect 16558 14384 16682 14426
rect 16390 14344 16392 14384
rect 16392 14344 16434 14384
rect 16434 14344 16474 14384
rect 16474 14344 16514 14384
rect 16558 14344 16598 14384
rect 16598 14344 16638 14384
rect 16638 14344 16680 14384
rect 16680 14344 16682 14384
rect 16390 14302 16514 14344
rect 16558 14302 16682 14344
rect 28390 14384 28514 14426
rect 28558 14384 28682 14426
rect 28390 14344 28392 14384
rect 28392 14344 28434 14384
rect 28434 14344 28474 14384
rect 28474 14344 28514 14384
rect 28558 14344 28598 14384
rect 28598 14344 28638 14384
rect 28638 14344 28680 14384
rect 28680 14344 28682 14384
rect 28390 14302 28514 14344
rect 28558 14302 28682 14344
rect 40390 14384 40514 14426
rect 40558 14384 40682 14426
rect 40390 14344 40392 14384
rect 40392 14344 40434 14384
rect 40434 14344 40474 14384
rect 40474 14344 40514 14384
rect 40558 14344 40598 14384
rect 40598 14344 40638 14384
rect 40638 14344 40680 14384
rect 40680 14344 40682 14384
rect 40390 14302 40514 14344
rect 40558 14302 40682 14344
rect 52390 14384 52514 14426
rect 52558 14384 52682 14426
rect 52390 14344 52392 14384
rect 52392 14344 52434 14384
rect 52434 14344 52474 14384
rect 52474 14344 52514 14384
rect 52558 14344 52598 14384
rect 52598 14344 52638 14384
rect 52638 14344 52680 14384
rect 52680 14344 52682 14384
rect 52390 14302 52514 14344
rect 52558 14302 52682 14344
rect 64390 14384 64514 14426
rect 64558 14384 64682 14426
rect 64390 14344 64392 14384
rect 64392 14344 64434 14384
rect 64434 14344 64474 14384
rect 64474 14344 64514 14384
rect 64558 14344 64598 14384
rect 64598 14344 64638 14384
rect 64638 14344 64680 14384
rect 64680 14344 64682 14384
rect 64390 14302 64514 14344
rect 64558 14302 64682 14344
rect 76390 14384 76514 14426
rect 76558 14384 76682 14426
rect 76390 14344 76392 14384
rect 76392 14344 76434 14384
rect 76434 14344 76474 14384
rect 76474 14344 76514 14384
rect 76558 14344 76598 14384
rect 76598 14344 76638 14384
rect 76638 14344 76680 14384
rect 76680 14344 76682 14384
rect 76390 14302 76514 14344
rect 76558 14302 76682 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 15150 13628 15274 13670
rect 15318 13628 15442 13670
rect 15150 13588 15152 13628
rect 15152 13588 15194 13628
rect 15194 13588 15234 13628
rect 15234 13588 15274 13628
rect 15318 13588 15358 13628
rect 15358 13588 15398 13628
rect 15398 13588 15440 13628
rect 15440 13588 15442 13628
rect 15150 13546 15274 13588
rect 15318 13546 15442 13588
rect 27150 13628 27274 13670
rect 27318 13628 27442 13670
rect 27150 13588 27152 13628
rect 27152 13588 27194 13628
rect 27194 13588 27234 13628
rect 27234 13588 27274 13628
rect 27318 13588 27358 13628
rect 27358 13588 27398 13628
rect 27398 13588 27440 13628
rect 27440 13588 27442 13628
rect 27150 13546 27274 13588
rect 27318 13546 27442 13588
rect 39150 13628 39274 13670
rect 39318 13628 39442 13670
rect 39150 13588 39152 13628
rect 39152 13588 39194 13628
rect 39194 13588 39234 13628
rect 39234 13588 39274 13628
rect 39318 13588 39358 13628
rect 39358 13588 39398 13628
rect 39398 13588 39440 13628
rect 39440 13588 39442 13628
rect 39150 13546 39274 13588
rect 39318 13546 39442 13588
rect 51150 13628 51274 13670
rect 51318 13628 51442 13670
rect 51150 13588 51152 13628
rect 51152 13588 51194 13628
rect 51194 13588 51234 13628
rect 51234 13588 51274 13628
rect 51318 13588 51358 13628
rect 51358 13588 51398 13628
rect 51398 13588 51440 13628
rect 51440 13588 51442 13628
rect 51150 13546 51274 13588
rect 51318 13546 51442 13588
rect 63150 13628 63274 13670
rect 63318 13628 63442 13670
rect 63150 13588 63152 13628
rect 63152 13588 63194 13628
rect 63194 13588 63234 13628
rect 63234 13588 63274 13628
rect 63318 13588 63358 13628
rect 63358 13588 63398 13628
rect 63398 13588 63440 13628
rect 63440 13588 63442 13628
rect 63150 13546 63274 13588
rect 63318 13546 63442 13588
rect 75150 13628 75274 13670
rect 75318 13628 75442 13670
rect 75150 13588 75152 13628
rect 75152 13588 75194 13628
rect 75194 13588 75234 13628
rect 75234 13588 75274 13628
rect 75318 13588 75358 13628
rect 75358 13588 75398 13628
rect 75398 13588 75440 13628
rect 75440 13588 75442 13628
rect 75150 13546 75274 13588
rect 75318 13546 75442 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 16390 12872 16514 12914
rect 16558 12872 16682 12914
rect 16390 12832 16392 12872
rect 16392 12832 16434 12872
rect 16434 12832 16474 12872
rect 16474 12832 16514 12872
rect 16558 12832 16598 12872
rect 16598 12832 16638 12872
rect 16638 12832 16680 12872
rect 16680 12832 16682 12872
rect 16390 12790 16514 12832
rect 16558 12790 16682 12832
rect 28390 12872 28514 12914
rect 28558 12872 28682 12914
rect 28390 12832 28392 12872
rect 28392 12832 28434 12872
rect 28434 12832 28474 12872
rect 28474 12832 28514 12872
rect 28558 12832 28598 12872
rect 28598 12832 28638 12872
rect 28638 12832 28680 12872
rect 28680 12832 28682 12872
rect 28390 12790 28514 12832
rect 28558 12790 28682 12832
rect 40390 12872 40514 12914
rect 40558 12872 40682 12914
rect 40390 12832 40392 12872
rect 40392 12832 40434 12872
rect 40434 12832 40474 12872
rect 40474 12832 40514 12872
rect 40558 12832 40598 12872
rect 40598 12832 40638 12872
rect 40638 12832 40680 12872
rect 40680 12832 40682 12872
rect 40390 12790 40514 12832
rect 40558 12790 40682 12832
rect 52390 12872 52514 12914
rect 52558 12872 52682 12914
rect 52390 12832 52392 12872
rect 52392 12832 52434 12872
rect 52434 12832 52474 12872
rect 52474 12832 52514 12872
rect 52558 12832 52598 12872
rect 52598 12832 52638 12872
rect 52638 12832 52680 12872
rect 52680 12832 52682 12872
rect 52390 12790 52514 12832
rect 52558 12790 52682 12832
rect 64390 12872 64514 12914
rect 64558 12872 64682 12914
rect 64390 12832 64392 12872
rect 64392 12832 64434 12872
rect 64434 12832 64474 12872
rect 64474 12832 64514 12872
rect 64558 12832 64598 12872
rect 64598 12832 64638 12872
rect 64638 12832 64680 12872
rect 64680 12832 64682 12872
rect 64390 12790 64514 12832
rect 64558 12790 64682 12832
rect 76390 12872 76514 12914
rect 76558 12872 76682 12914
rect 76390 12832 76392 12872
rect 76392 12832 76434 12872
rect 76434 12832 76474 12872
rect 76474 12832 76514 12872
rect 76558 12832 76598 12872
rect 76598 12832 76638 12872
rect 76638 12832 76680 12872
rect 76680 12832 76682 12872
rect 76390 12790 76514 12832
rect 76558 12790 76682 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 15150 12116 15274 12158
rect 15318 12116 15442 12158
rect 15150 12076 15152 12116
rect 15152 12076 15194 12116
rect 15194 12076 15234 12116
rect 15234 12076 15274 12116
rect 15318 12076 15358 12116
rect 15358 12076 15398 12116
rect 15398 12076 15440 12116
rect 15440 12076 15442 12116
rect 15150 12034 15274 12076
rect 15318 12034 15442 12076
rect 27150 12116 27274 12158
rect 27318 12116 27442 12158
rect 27150 12076 27152 12116
rect 27152 12076 27194 12116
rect 27194 12076 27234 12116
rect 27234 12076 27274 12116
rect 27318 12076 27358 12116
rect 27358 12076 27398 12116
rect 27398 12076 27440 12116
rect 27440 12076 27442 12116
rect 27150 12034 27274 12076
rect 27318 12034 27442 12076
rect 39150 12116 39274 12158
rect 39318 12116 39442 12158
rect 39150 12076 39152 12116
rect 39152 12076 39194 12116
rect 39194 12076 39234 12116
rect 39234 12076 39274 12116
rect 39318 12076 39358 12116
rect 39358 12076 39398 12116
rect 39398 12076 39440 12116
rect 39440 12076 39442 12116
rect 39150 12034 39274 12076
rect 39318 12034 39442 12076
rect 51150 12116 51274 12158
rect 51318 12116 51442 12158
rect 51150 12076 51152 12116
rect 51152 12076 51194 12116
rect 51194 12076 51234 12116
rect 51234 12076 51274 12116
rect 51318 12076 51358 12116
rect 51358 12076 51398 12116
rect 51398 12076 51440 12116
rect 51440 12076 51442 12116
rect 51150 12034 51274 12076
rect 51318 12034 51442 12076
rect 63150 12116 63274 12158
rect 63318 12116 63442 12158
rect 63150 12076 63152 12116
rect 63152 12076 63194 12116
rect 63194 12076 63234 12116
rect 63234 12076 63274 12116
rect 63318 12076 63358 12116
rect 63358 12076 63398 12116
rect 63398 12076 63440 12116
rect 63440 12076 63442 12116
rect 63150 12034 63274 12076
rect 63318 12034 63442 12076
rect 75150 12116 75274 12158
rect 75318 12116 75442 12158
rect 75150 12076 75152 12116
rect 75152 12076 75194 12116
rect 75194 12076 75234 12116
rect 75234 12076 75274 12116
rect 75318 12076 75358 12116
rect 75358 12076 75398 12116
rect 75398 12076 75440 12116
rect 75440 12076 75442 12116
rect 75150 12034 75274 12076
rect 75318 12034 75442 12076
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 16390 11360 16514 11402
rect 16558 11360 16682 11402
rect 16390 11320 16392 11360
rect 16392 11320 16434 11360
rect 16434 11320 16474 11360
rect 16474 11320 16514 11360
rect 16558 11320 16598 11360
rect 16598 11320 16638 11360
rect 16638 11320 16680 11360
rect 16680 11320 16682 11360
rect 16390 11278 16514 11320
rect 16558 11278 16682 11320
rect 28390 11360 28514 11402
rect 28558 11360 28682 11402
rect 28390 11320 28392 11360
rect 28392 11320 28434 11360
rect 28434 11320 28474 11360
rect 28474 11320 28514 11360
rect 28558 11320 28598 11360
rect 28598 11320 28638 11360
rect 28638 11320 28680 11360
rect 28680 11320 28682 11360
rect 28390 11278 28514 11320
rect 28558 11278 28682 11320
rect 40390 11360 40514 11402
rect 40558 11360 40682 11402
rect 40390 11320 40392 11360
rect 40392 11320 40434 11360
rect 40434 11320 40474 11360
rect 40474 11320 40514 11360
rect 40558 11320 40598 11360
rect 40598 11320 40638 11360
rect 40638 11320 40680 11360
rect 40680 11320 40682 11360
rect 40390 11278 40514 11320
rect 40558 11278 40682 11320
rect 52390 11360 52514 11402
rect 52558 11360 52682 11402
rect 52390 11320 52392 11360
rect 52392 11320 52434 11360
rect 52434 11320 52474 11360
rect 52474 11320 52514 11360
rect 52558 11320 52598 11360
rect 52598 11320 52638 11360
rect 52638 11320 52680 11360
rect 52680 11320 52682 11360
rect 52390 11278 52514 11320
rect 52558 11278 52682 11320
rect 64390 11360 64514 11402
rect 64558 11360 64682 11402
rect 64390 11320 64392 11360
rect 64392 11320 64434 11360
rect 64434 11320 64474 11360
rect 64474 11320 64514 11360
rect 64558 11320 64598 11360
rect 64598 11320 64638 11360
rect 64638 11320 64680 11360
rect 64680 11320 64682 11360
rect 64390 11278 64514 11320
rect 64558 11278 64682 11320
rect 76390 11360 76514 11402
rect 76558 11360 76682 11402
rect 76390 11320 76392 11360
rect 76392 11320 76434 11360
rect 76434 11320 76474 11360
rect 76474 11320 76514 11360
rect 76558 11320 76598 11360
rect 76598 11320 76638 11360
rect 76638 11320 76680 11360
rect 76680 11320 76682 11360
rect 76390 11278 76514 11320
rect 76558 11278 76682 11320
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 15150 10604 15274 10646
rect 15318 10604 15442 10646
rect 15150 10564 15152 10604
rect 15152 10564 15194 10604
rect 15194 10564 15234 10604
rect 15234 10564 15274 10604
rect 15318 10564 15358 10604
rect 15358 10564 15398 10604
rect 15398 10564 15440 10604
rect 15440 10564 15442 10604
rect 15150 10522 15274 10564
rect 15318 10522 15442 10564
rect 27150 10604 27274 10646
rect 27318 10604 27442 10646
rect 27150 10564 27152 10604
rect 27152 10564 27194 10604
rect 27194 10564 27234 10604
rect 27234 10564 27274 10604
rect 27318 10564 27358 10604
rect 27358 10564 27398 10604
rect 27398 10564 27440 10604
rect 27440 10564 27442 10604
rect 27150 10522 27274 10564
rect 27318 10522 27442 10564
rect 39150 10604 39274 10646
rect 39318 10604 39442 10646
rect 39150 10564 39152 10604
rect 39152 10564 39194 10604
rect 39194 10564 39234 10604
rect 39234 10564 39274 10604
rect 39318 10564 39358 10604
rect 39358 10564 39398 10604
rect 39398 10564 39440 10604
rect 39440 10564 39442 10604
rect 39150 10522 39274 10564
rect 39318 10522 39442 10564
rect 51150 10604 51274 10646
rect 51318 10604 51442 10646
rect 51150 10564 51152 10604
rect 51152 10564 51194 10604
rect 51194 10564 51234 10604
rect 51234 10564 51274 10604
rect 51318 10564 51358 10604
rect 51358 10564 51398 10604
rect 51398 10564 51440 10604
rect 51440 10564 51442 10604
rect 51150 10522 51274 10564
rect 51318 10522 51442 10564
rect 63150 10604 63274 10646
rect 63318 10604 63442 10646
rect 63150 10564 63152 10604
rect 63152 10564 63194 10604
rect 63194 10564 63234 10604
rect 63234 10564 63274 10604
rect 63318 10564 63358 10604
rect 63358 10564 63398 10604
rect 63398 10564 63440 10604
rect 63440 10564 63442 10604
rect 63150 10522 63274 10564
rect 63318 10522 63442 10564
rect 75150 10604 75274 10646
rect 75318 10604 75442 10646
rect 75150 10564 75152 10604
rect 75152 10564 75194 10604
rect 75194 10564 75234 10604
rect 75234 10564 75274 10604
rect 75318 10564 75358 10604
rect 75358 10564 75398 10604
rect 75398 10564 75440 10604
rect 75440 10564 75442 10604
rect 75150 10522 75274 10564
rect 75318 10522 75442 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 16390 9848 16514 9890
rect 16558 9848 16682 9890
rect 16390 9808 16392 9848
rect 16392 9808 16434 9848
rect 16434 9808 16474 9848
rect 16474 9808 16514 9848
rect 16558 9808 16598 9848
rect 16598 9808 16638 9848
rect 16638 9808 16680 9848
rect 16680 9808 16682 9848
rect 16390 9766 16514 9808
rect 16558 9766 16682 9808
rect 28390 9848 28514 9890
rect 28558 9848 28682 9890
rect 28390 9808 28392 9848
rect 28392 9808 28434 9848
rect 28434 9808 28474 9848
rect 28474 9808 28514 9848
rect 28558 9808 28598 9848
rect 28598 9808 28638 9848
rect 28638 9808 28680 9848
rect 28680 9808 28682 9848
rect 28390 9766 28514 9808
rect 28558 9766 28682 9808
rect 40390 9848 40514 9890
rect 40558 9848 40682 9890
rect 40390 9808 40392 9848
rect 40392 9808 40434 9848
rect 40434 9808 40474 9848
rect 40474 9808 40514 9848
rect 40558 9808 40598 9848
rect 40598 9808 40638 9848
rect 40638 9808 40680 9848
rect 40680 9808 40682 9848
rect 40390 9766 40514 9808
rect 40558 9766 40682 9808
rect 52390 9848 52514 9890
rect 52558 9848 52682 9890
rect 52390 9808 52392 9848
rect 52392 9808 52434 9848
rect 52434 9808 52474 9848
rect 52474 9808 52514 9848
rect 52558 9808 52598 9848
rect 52598 9808 52638 9848
rect 52638 9808 52680 9848
rect 52680 9808 52682 9848
rect 52390 9766 52514 9808
rect 52558 9766 52682 9808
rect 64390 9848 64514 9890
rect 64558 9848 64682 9890
rect 64390 9808 64392 9848
rect 64392 9808 64434 9848
rect 64434 9808 64474 9848
rect 64474 9808 64514 9848
rect 64558 9808 64598 9848
rect 64598 9808 64638 9848
rect 64638 9808 64680 9848
rect 64680 9808 64682 9848
rect 64390 9766 64514 9808
rect 64558 9766 64682 9808
rect 76390 9848 76514 9890
rect 76558 9848 76682 9890
rect 76390 9808 76392 9848
rect 76392 9808 76434 9848
rect 76434 9808 76474 9848
rect 76474 9808 76514 9848
rect 76558 9808 76598 9848
rect 76598 9808 76638 9848
rect 76638 9808 76680 9848
rect 76680 9808 76682 9848
rect 76390 9766 76514 9808
rect 76558 9766 76682 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 15150 9092 15274 9134
rect 15318 9092 15442 9134
rect 15150 9052 15152 9092
rect 15152 9052 15194 9092
rect 15194 9052 15234 9092
rect 15234 9052 15274 9092
rect 15318 9052 15358 9092
rect 15358 9052 15398 9092
rect 15398 9052 15440 9092
rect 15440 9052 15442 9092
rect 15150 9010 15274 9052
rect 15318 9010 15442 9052
rect 27150 9092 27274 9134
rect 27318 9092 27442 9134
rect 27150 9052 27152 9092
rect 27152 9052 27194 9092
rect 27194 9052 27234 9092
rect 27234 9052 27274 9092
rect 27318 9052 27358 9092
rect 27358 9052 27398 9092
rect 27398 9052 27440 9092
rect 27440 9052 27442 9092
rect 27150 9010 27274 9052
rect 27318 9010 27442 9052
rect 39150 9092 39274 9134
rect 39318 9092 39442 9134
rect 39150 9052 39152 9092
rect 39152 9052 39194 9092
rect 39194 9052 39234 9092
rect 39234 9052 39274 9092
rect 39318 9052 39358 9092
rect 39358 9052 39398 9092
rect 39398 9052 39440 9092
rect 39440 9052 39442 9092
rect 39150 9010 39274 9052
rect 39318 9010 39442 9052
rect 51150 9092 51274 9134
rect 51318 9092 51442 9134
rect 51150 9052 51152 9092
rect 51152 9052 51194 9092
rect 51194 9052 51234 9092
rect 51234 9052 51274 9092
rect 51318 9052 51358 9092
rect 51358 9052 51398 9092
rect 51398 9052 51440 9092
rect 51440 9052 51442 9092
rect 51150 9010 51274 9052
rect 51318 9010 51442 9052
rect 63150 9092 63274 9134
rect 63318 9092 63442 9134
rect 63150 9052 63152 9092
rect 63152 9052 63194 9092
rect 63194 9052 63234 9092
rect 63234 9052 63274 9092
rect 63318 9052 63358 9092
rect 63358 9052 63398 9092
rect 63398 9052 63440 9092
rect 63440 9052 63442 9092
rect 63150 9010 63274 9052
rect 63318 9010 63442 9052
rect 75150 9092 75274 9134
rect 75318 9092 75442 9134
rect 75150 9052 75152 9092
rect 75152 9052 75194 9092
rect 75194 9052 75234 9092
rect 75234 9052 75274 9092
rect 75318 9052 75358 9092
rect 75358 9052 75398 9092
rect 75398 9052 75440 9092
rect 75440 9052 75442 9092
rect 75150 9010 75274 9052
rect 75318 9010 75442 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 16390 8336 16514 8378
rect 16558 8336 16682 8378
rect 16390 8296 16392 8336
rect 16392 8296 16434 8336
rect 16434 8296 16474 8336
rect 16474 8296 16514 8336
rect 16558 8296 16598 8336
rect 16598 8296 16638 8336
rect 16638 8296 16680 8336
rect 16680 8296 16682 8336
rect 16390 8254 16514 8296
rect 16558 8254 16682 8296
rect 28390 8336 28514 8378
rect 28558 8336 28682 8378
rect 28390 8296 28392 8336
rect 28392 8296 28434 8336
rect 28434 8296 28474 8336
rect 28474 8296 28514 8336
rect 28558 8296 28598 8336
rect 28598 8296 28638 8336
rect 28638 8296 28680 8336
rect 28680 8296 28682 8336
rect 28390 8254 28514 8296
rect 28558 8254 28682 8296
rect 40390 8336 40514 8378
rect 40558 8336 40682 8378
rect 40390 8296 40392 8336
rect 40392 8296 40434 8336
rect 40434 8296 40474 8336
rect 40474 8296 40514 8336
rect 40558 8296 40598 8336
rect 40598 8296 40638 8336
rect 40638 8296 40680 8336
rect 40680 8296 40682 8336
rect 40390 8254 40514 8296
rect 40558 8254 40682 8296
rect 52390 8336 52514 8378
rect 52558 8336 52682 8378
rect 52390 8296 52392 8336
rect 52392 8296 52434 8336
rect 52434 8296 52474 8336
rect 52474 8296 52514 8336
rect 52558 8296 52598 8336
rect 52598 8296 52638 8336
rect 52638 8296 52680 8336
rect 52680 8296 52682 8336
rect 52390 8254 52514 8296
rect 52558 8254 52682 8296
rect 64390 8336 64514 8378
rect 64558 8336 64682 8378
rect 64390 8296 64392 8336
rect 64392 8296 64434 8336
rect 64434 8296 64474 8336
rect 64474 8296 64514 8336
rect 64558 8296 64598 8336
rect 64598 8296 64638 8336
rect 64638 8296 64680 8336
rect 64680 8296 64682 8336
rect 64390 8254 64514 8296
rect 64558 8254 64682 8296
rect 76390 8336 76514 8378
rect 76558 8336 76682 8378
rect 76390 8296 76392 8336
rect 76392 8296 76434 8336
rect 76434 8296 76474 8336
rect 76474 8296 76514 8336
rect 76558 8296 76598 8336
rect 76598 8296 76638 8336
rect 76638 8296 76680 8336
rect 76680 8296 76682 8336
rect 76390 8254 76514 8296
rect 76558 8254 76682 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 15150 7580 15274 7622
rect 15318 7580 15442 7622
rect 15150 7540 15152 7580
rect 15152 7540 15194 7580
rect 15194 7540 15234 7580
rect 15234 7540 15274 7580
rect 15318 7540 15358 7580
rect 15358 7540 15398 7580
rect 15398 7540 15440 7580
rect 15440 7540 15442 7580
rect 15150 7498 15274 7540
rect 15318 7498 15442 7540
rect 27150 7580 27274 7622
rect 27318 7580 27442 7622
rect 27150 7540 27152 7580
rect 27152 7540 27194 7580
rect 27194 7540 27234 7580
rect 27234 7540 27274 7580
rect 27318 7540 27358 7580
rect 27358 7540 27398 7580
rect 27398 7540 27440 7580
rect 27440 7540 27442 7580
rect 27150 7498 27274 7540
rect 27318 7498 27442 7540
rect 39150 7580 39274 7622
rect 39318 7580 39442 7622
rect 39150 7540 39152 7580
rect 39152 7540 39194 7580
rect 39194 7540 39234 7580
rect 39234 7540 39274 7580
rect 39318 7540 39358 7580
rect 39358 7540 39398 7580
rect 39398 7540 39440 7580
rect 39440 7540 39442 7580
rect 39150 7498 39274 7540
rect 39318 7498 39442 7540
rect 51150 7580 51274 7622
rect 51318 7580 51442 7622
rect 51150 7540 51152 7580
rect 51152 7540 51194 7580
rect 51194 7540 51234 7580
rect 51234 7540 51274 7580
rect 51318 7540 51358 7580
rect 51358 7540 51398 7580
rect 51398 7540 51440 7580
rect 51440 7540 51442 7580
rect 51150 7498 51274 7540
rect 51318 7498 51442 7540
rect 63150 7580 63274 7622
rect 63318 7580 63442 7622
rect 63150 7540 63152 7580
rect 63152 7540 63194 7580
rect 63194 7540 63234 7580
rect 63234 7540 63274 7580
rect 63318 7540 63358 7580
rect 63358 7540 63398 7580
rect 63398 7540 63440 7580
rect 63440 7540 63442 7580
rect 63150 7498 63274 7540
rect 63318 7498 63442 7540
rect 75150 7580 75274 7622
rect 75318 7580 75442 7622
rect 75150 7540 75152 7580
rect 75152 7540 75194 7580
rect 75194 7540 75234 7580
rect 75234 7540 75274 7580
rect 75318 7540 75358 7580
rect 75358 7540 75398 7580
rect 75398 7540 75440 7580
rect 75440 7540 75442 7580
rect 75150 7498 75274 7540
rect 75318 7498 75442 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 16390 6824 16514 6866
rect 16558 6824 16682 6866
rect 16390 6784 16392 6824
rect 16392 6784 16434 6824
rect 16434 6784 16474 6824
rect 16474 6784 16514 6824
rect 16558 6784 16598 6824
rect 16598 6784 16638 6824
rect 16638 6784 16680 6824
rect 16680 6784 16682 6824
rect 16390 6742 16514 6784
rect 16558 6742 16682 6784
rect 28390 6824 28514 6866
rect 28558 6824 28682 6866
rect 28390 6784 28392 6824
rect 28392 6784 28434 6824
rect 28434 6784 28474 6824
rect 28474 6784 28514 6824
rect 28558 6784 28598 6824
rect 28598 6784 28638 6824
rect 28638 6784 28680 6824
rect 28680 6784 28682 6824
rect 28390 6742 28514 6784
rect 28558 6742 28682 6784
rect 40390 6824 40514 6866
rect 40558 6824 40682 6866
rect 40390 6784 40392 6824
rect 40392 6784 40434 6824
rect 40434 6784 40474 6824
rect 40474 6784 40514 6824
rect 40558 6784 40598 6824
rect 40598 6784 40638 6824
rect 40638 6784 40680 6824
rect 40680 6784 40682 6824
rect 40390 6742 40514 6784
rect 40558 6742 40682 6784
rect 52390 6824 52514 6866
rect 52558 6824 52682 6866
rect 52390 6784 52392 6824
rect 52392 6784 52434 6824
rect 52434 6784 52474 6824
rect 52474 6784 52514 6824
rect 52558 6784 52598 6824
rect 52598 6784 52638 6824
rect 52638 6784 52680 6824
rect 52680 6784 52682 6824
rect 52390 6742 52514 6784
rect 52558 6742 52682 6784
rect 64390 6824 64514 6866
rect 64558 6824 64682 6866
rect 64390 6784 64392 6824
rect 64392 6784 64434 6824
rect 64434 6784 64474 6824
rect 64474 6784 64514 6824
rect 64558 6784 64598 6824
rect 64598 6784 64638 6824
rect 64638 6784 64680 6824
rect 64680 6784 64682 6824
rect 64390 6742 64514 6784
rect 64558 6742 64682 6784
rect 76390 6824 76514 6866
rect 76558 6824 76682 6866
rect 76390 6784 76392 6824
rect 76392 6784 76434 6824
rect 76434 6784 76474 6824
rect 76474 6784 76514 6824
rect 76558 6784 76598 6824
rect 76598 6784 76638 6824
rect 76638 6784 76680 6824
rect 76680 6784 76682 6824
rect 76390 6742 76514 6784
rect 76558 6742 76682 6784
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 15150 6068 15274 6110
rect 15318 6068 15442 6110
rect 15150 6028 15152 6068
rect 15152 6028 15194 6068
rect 15194 6028 15234 6068
rect 15234 6028 15274 6068
rect 15318 6028 15358 6068
rect 15358 6028 15398 6068
rect 15398 6028 15440 6068
rect 15440 6028 15442 6068
rect 15150 5986 15274 6028
rect 15318 5986 15442 6028
rect 27150 6068 27274 6110
rect 27318 6068 27442 6110
rect 27150 6028 27152 6068
rect 27152 6028 27194 6068
rect 27194 6028 27234 6068
rect 27234 6028 27274 6068
rect 27318 6028 27358 6068
rect 27358 6028 27398 6068
rect 27398 6028 27440 6068
rect 27440 6028 27442 6068
rect 27150 5986 27274 6028
rect 27318 5986 27442 6028
rect 39150 6068 39274 6110
rect 39318 6068 39442 6110
rect 39150 6028 39152 6068
rect 39152 6028 39194 6068
rect 39194 6028 39234 6068
rect 39234 6028 39274 6068
rect 39318 6028 39358 6068
rect 39358 6028 39398 6068
rect 39398 6028 39440 6068
rect 39440 6028 39442 6068
rect 39150 5986 39274 6028
rect 39318 5986 39442 6028
rect 51150 6068 51274 6110
rect 51318 6068 51442 6110
rect 51150 6028 51152 6068
rect 51152 6028 51194 6068
rect 51194 6028 51234 6068
rect 51234 6028 51274 6068
rect 51318 6028 51358 6068
rect 51358 6028 51398 6068
rect 51398 6028 51440 6068
rect 51440 6028 51442 6068
rect 51150 5986 51274 6028
rect 51318 5986 51442 6028
rect 63150 6068 63274 6110
rect 63318 6068 63442 6110
rect 63150 6028 63152 6068
rect 63152 6028 63194 6068
rect 63194 6028 63234 6068
rect 63234 6028 63274 6068
rect 63318 6028 63358 6068
rect 63358 6028 63398 6068
rect 63398 6028 63440 6068
rect 63440 6028 63442 6068
rect 63150 5986 63274 6028
rect 63318 5986 63442 6028
rect 75150 6068 75274 6110
rect 75318 6068 75442 6110
rect 75150 6028 75152 6068
rect 75152 6028 75194 6068
rect 75194 6028 75234 6068
rect 75234 6028 75274 6068
rect 75318 6028 75358 6068
rect 75358 6028 75398 6068
rect 75398 6028 75440 6068
rect 75440 6028 75442 6068
rect 75150 5986 75274 6028
rect 75318 5986 75442 6028
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 16390 5312 16514 5354
rect 16558 5312 16682 5354
rect 16390 5272 16392 5312
rect 16392 5272 16434 5312
rect 16434 5272 16474 5312
rect 16474 5272 16514 5312
rect 16558 5272 16598 5312
rect 16598 5272 16638 5312
rect 16638 5272 16680 5312
rect 16680 5272 16682 5312
rect 16390 5230 16514 5272
rect 16558 5230 16682 5272
rect 28390 5312 28514 5354
rect 28558 5312 28682 5354
rect 28390 5272 28392 5312
rect 28392 5272 28434 5312
rect 28434 5272 28474 5312
rect 28474 5272 28514 5312
rect 28558 5272 28598 5312
rect 28598 5272 28638 5312
rect 28638 5272 28680 5312
rect 28680 5272 28682 5312
rect 28390 5230 28514 5272
rect 28558 5230 28682 5272
rect 40390 5312 40514 5354
rect 40558 5312 40682 5354
rect 40390 5272 40392 5312
rect 40392 5272 40434 5312
rect 40434 5272 40474 5312
rect 40474 5272 40514 5312
rect 40558 5272 40598 5312
rect 40598 5272 40638 5312
rect 40638 5272 40680 5312
rect 40680 5272 40682 5312
rect 40390 5230 40514 5272
rect 40558 5230 40682 5272
rect 52390 5312 52514 5354
rect 52558 5312 52682 5354
rect 52390 5272 52392 5312
rect 52392 5272 52434 5312
rect 52434 5272 52474 5312
rect 52474 5272 52514 5312
rect 52558 5272 52598 5312
rect 52598 5272 52638 5312
rect 52638 5272 52680 5312
rect 52680 5272 52682 5312
rect 52390 5230 52514 5272
rect 52558 5230 52682 5272
rect 64390 5312 64514 5354
rect 64558 5312 64682 5354
rect 64390 5272 64392 5312
rect 64392 5272 64434 5312
rect 64434 5272 64474 5312
rect 64474 5272 64514 5312
rect 64558 5272 64598 5312
rect 64598 5272 64638 5312
rect 64638 5272 64680 5312
rect 64680 5272 64682 5312
rect 64390 5230 64514 5272
rect 64558 5230 64682 5272
rect 76390 5312 76514 5354
rect 76558 5312 76682 5354
rect 76390 5272 76392 5312
rect 76392 5272 76434 5312
rect 76434 5272 76474 5312
rect 76474 5272 76514 5312
rect 76558 5272 76598 5312
rect 76598 5272 76638 5312
rect 76638 5272 76680 5312
rect 76680 5272 76682 5312
rect 76390 5230 76514 5272
rect 76558 5230 76682 5272
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 15150 4556 15274 4598
rect 15318 4556 15442 4598
rect 15150 4516 15152 4556
rect 15152 4516 15194 4556
rect 15194 4516 15234 4556
rect 15234 4516 15274 4556
rect 15318 4516 15358 4556
rect 15358 4516 15398 4556
rect 15398 4516 15440 4556
rect 15440 4516 15442 4556
rect 15150 4474 15274 4516
rect 15318 4474 15442 4516
rect 27150 4556 27274 4598
rect 27318 4556 27442 4598
rect 27150 4516 27152 4556
rect 27152 4516 27194 4556
rect 27194 4516 27234 4556
rect 27234 4516 27274 4556
rect 27318 4516 27358 4556
rect 27358 4516 27398 4556
rect 27398 4516 27440 4556
rect 27440 4516 27442 4556
rect 27150 4474 27274 4516
rect 27318 4474 27442 4516
rect 39150 4556 39274 4598
rect 39318 4556 39442 4598
rect 39150 4516 39152 4556
rect 39152 4516 39194 4556
rect 39194 4516 39234 4556
rect 39234 4516 39274 4556
rect 39318 4516 39358 4556
rect 39358 4516 39398 4556
rect 39398 4516 39440 4556
rect 39440 4516 39442 4556
rect 39150 4474 39274 4516
rect 39318 4474 39442 4516
rect 51150 4556 51274 4598
rect 51318 4556 51442 4598
rect 51150 4516 51152 4556
rect 51152 4516 51194 4556
rect 51194 4516 51234 4556
rect 51234 4516 51274 4556
rect 51318 4516 51358 4556
rect 51358 4516 51398 4556
rect 51398 4516 51440 4556
rect 51440 4516 51442 4556
rect 51150 4474 51274 4516
rect 51318 4474 51442 4516
rect 63150 4556 63274 4598
rect 63318 4556 63442 4598
rect 63150 4516 63152 4556
rect 63152 4516 63194 4556
rect 63194 4516 63234 4556
rect 63234 4516 63274 4556
rect 63318 4516 63358 4556
rect 63358 4516 63398 4556
rect 63398 4516 63440 4556
rect 63440 4516 63442 4556
rect 63150 4474 63274 4516
rect 63318 4474 63442 4516
rect 75150 4556 75274 4598
rect 75318 4556 75442 4598
rect 75150 4516 75152 4556
rect 75152 4516 75194 4556
rect 75194 4516 75234 4556
rect 75234 4516 75274 4556
rect 75318 4516 75358 4556
rect 75358 4516 75398 4556
rect 75398 4516 75440 4556
rect 75440 4516 75442 4556
rect 75150 4474 75274 4516
rect 75318 4474 75442 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 16390 3800 16514 3842
rect 16558 3800 16682 3842
rect 16390 3760 16392 3800
rect 16392 3760 16434 3800
rect 16434 3760 16474 3800
rect 16474 3760 16514 3800
rect 16558 3760 16598 3800
rect 16598 3760 16638 3800
rect 16638 3760 16680 3800
rect 16680 3760 16682 3800
rect 16390 3718 16514 3760
rect 16558 3718 16682 3760
rect 28390 3800 28514 3842
rect 28558 3800 28682 3842
rect 28390 3760 28392 3800
rect 28392 3760 28434 3800
rect 28434 3760 28474 3800
rect 28474 3760 28514 3800
rect 28558 3760 28598 3800
rect 28598 3760 28638 3800
rect 28638 3760 28680 3800
rect 28680 3760 28682 3800
rect 28390 3718 28514 3760
rect 28558 3718 28682 3760
rect 40390 3800 40514 3842
rect 40558 3800 40682 3842
rect 40390 3760 40392 3800
rect 40392 3760 40434 3800
rect 40434 3760 40474 3800
rect 40474 3760 40514 3800
rect 40558 3760 40598 3800
rect 40598 3760 40638 3800
rect 40638 3760 40680 3800
rect 40680 3760 40682 3800
rect 40390 3718 40514 3760
rect 40558 3718 40682 3760
rect 52390 3800 52514 3842
rect 52558 3800 52682 3842
rect 52390 3760 52392 3800
rect 52392 3760 52434 3800
rect 52434 3760 52474 3800
rect 52474 3760 52514 3800
rect 52558 3760 52598 3800
rect 52598 3760 52638 3800
rect 52638 3760 52680 3800
rect 52680 3760 52682 3800
rect 52390 3718 52514 3760
rect 52558 3718 52682 3760
rect 64390 3800 64514 3842
rect 64558 3800 64682 3842
rect 64390 3760 64392 3800
rect 64392 3760 64434 3800
rect 64434 3760 64474 3800
rect 64474 3760 64514 3800
rect 64558 3760 64598 3800
rect 64598 3760 64638 3800
rect 64638 3760 64680 3800
rect 64680 3760 64682 3800
rect 64390 3718 64514 3760
rect 64558 3718 64682 3760
rect 76390 3800 76514 3842
rect 76558 3800 76682 3842
rect 76390 3760 76392 3800
rect 76392 3760 76434 3800
rect 76434 3760 76474 3800
rect 76474 3760 76514 3800
rect 76558 3760 76598 3800
rect 76598 3760 76638 3800
rect 76638 3760 76680 3800
rect 76680 3760 76682 3800
rect 76390 3718 76514 3760
rect 76558 3718 76682 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 15150 3044 15274 3086
rect 15318 3044 15442 3086
rect 15150 3004 15152 3044
rect 15152 3004 15194 3044
rect 15194 3004 15234 3044
rect 15234 3004 15274 3044
rect 15318 3004 15358 3044
rect 15358 3004 15398 3044
rect 15398 3004 15440 3044
rect 15440 3004 15442 3044
rect 15150 2962 15274 3004
rect 15318 2962 15442 3004
rect 27150 3044 27274 3086
rect 27318 3044 27442 3086
rect 27150 3004 27152 3044
rect 27152 3004 27194 3044
rect 27194 3004 27234 3044
rect 27234 3004 27274 3044
rect 27318 3004 27358 3044
rect 27358 3004 27398 3044
rect 27398 3004 27440 3044
rect 27440 3004 27442 3044
rect 27150 2962 27274 3004
rect 27318 2962 27442 3004
rect 39150 3044 39274 3086
rect 39318 3044 39442 3086
rect 39150 3004 39152 3044
rect 39152 3004 39194 3044
rect 39194 3004 39234 3044
rect 39234 3004 39274 3044
rect 39318 3004 39358 3044
rect 39358 3004 39398 3044
rect 39398 3004 39440 3044
rect 39440 3004 39442 3044
rect 39150 2962 39274 3004
rect 39318 2962 39442 3004
rect 51150 3044 51274 3086
rect 51318 3044 51442 3086
rect 51150 3004 51152 3044
rect 51152 3004 51194 3044
rect 51194 3004 51234 3044
rect 51234 3004 51274 3044
rect 51318 3004 51358 3044
rect 51358 3004 51398 3044
rect 51398 3004 51440 3044
rect 51440 3004 51442 3044
rect 51150 2962 51274 3004
rect 51318 2962 51442 3004
rect 63150 3044 63274 3086
rect 63318 3044 63442 3086
rect 63150 3004 63152 3044
rect 63152 3004 63194 3044
rect 63194 3004 63234 3044
rect 63234 3004 63274 3044
rect 63318 3004 63358 3044
rect 63358 3004 63398 3044
rect 63398 3004 63440 3044
rect 63440 3004 63442 3044
rect 63150 2962 63274 3004
rect 63318 2962 63442 3004
rect 75150 3044 75274 3086
rect 75318 3044 75442 3086
rect 75150 3004 75152 3044
rect 75152 3004 75194 3044
rect 75194 3004 75234 3044
rect 75234 3004 75274 3044
rect 75318 3004 75358 3044
rect 75358 3004 75398 3044
rect 75398 3004 75440 3044
rect 75440 3004 75442 3044
rect 75150 2962 75274 3004
rect 75318 2962 75442 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 16390 2288 16514 2330
rect 16558 2288 16682 2330
rect 16390 2248 16392 2288
rect 16392 2248 16434 2288
rect 16434 2248 16474 2288
rect 16474 2248 16514 2288
rect 16558 2248 16598 2288
rect 16598 2248 16638 2288
rect 16638 2248 16680 2288
rect 16680 2248 16682 2288
rect 16390 2206 16514 2248
rect 16558 2206 16682 2248
rect 28390 2288 28514 2330
rect 28558 2288 28682 2330
rect 28390 2248 28392 2288
rect 28392 2248 28434 2288
rect 28434 2248 28474 2288
rect 28474 2248 28514 2288
rect 28558 2248 28598 2288
rect 28598 2248 28638 2288
rect 28638 2248 28680 2288
rect 28680 2248 28682 2288
rect 28390 2206 28514 2248
rect 28558 2206 28682 2248
rect 40390 2288 40514 2330
rect 40558 2288 40682 2330
rect 40390 2248 40392 2288
rect 40392 2248 40434 2288
rect 40434 2248 40474 2288
rect 40474 2248 40514 2288
rect 40558 2248 40598 2288
rect 40598 2248 40638 2288
rect 40638 2248 40680 2288
rect 40680 2248 40682 2288
rect 40390 2206 40514 2248
rect 40558 2206 40682 2248
rect 52390 2288 52514 2330
rect 52558 2288 52682 2330
rect 52390 2248 52392 2288
rect 52392 2248 52434 2288
rect 52434 2248 52474 2288
rect 52474 2248 52514 2288
rect 52558 2248 52598 2288
rect 52598 2248 52638 2288
rect 52638 2248 52680 2288
rect 52680 2248 52682 2288
rect 52390 2206 52514 2248
rect 52558 2206 52682 2248
rect 64390 2288 64514 2330
rect 64558 2288 64682 2330
rect 64390 2248 64392 2288
rect 64392 2248 64434 2288
rect 64434 2248 64474 2288
rect 64474 2248 64514 2288
rect 64558 2248 64598 2288
rect 64598 2248 64638 2288
rect 64638 2248 64680 2288
rect 64680 2248 64682 2288
rect 64390 2206 64514 2248
rect 64558 2206 64682 2248
rect 76390 2288 76514 2330
rect 76558 2288 76682 2330
rect 76390 2248 76392 2288
rect 76392 2248 76434 2288
rect 76434 2248 76474 2288
rect 76474 2248 76514 2288
rect 76558 2248 76598 2288
rect 76598 2248 76638 2288
rect 76638 2248 76680 2288
rect 76680 2248 76682 2288
rect 76390 2206 76514 2248
rect 76558 2206 76682 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 15150 1532 15274 1574
rect 15318 1532 15442 1574
rect 15150 1492 15152 1532
rect 15152 1492 15194 1532
rect 15194 1492 15234 1532
rect 15234 1492 15274 1532
rect 15318 1492 15358 1532
rect 15358 1492 15398 1532
rect 15398 1492 15440 1532
rect 15440 1492 15442 1532
rect 15150 1450 15274 1492
rect 15318 1450 15442 1492
rect 27150 1532 27274 1574
rect 27318 1532 27442 1574
rect 27150 1492 27152 1532
rect 27152 1492 27194 1532
rect 27194 1492 27234 1532
rect 27234 1492 27274 1532
rect 27318 1492 27358 1532
rect 27358 1492 27398 1532
rect 27398 1492 27440 1532
rect 27440 1492 27442 1532
rect 27150 1450 27274 1492
rect 27318 1450 27442 1492
rect 39150 1532 39274 1574
rect 39318 1532 39442 1574
rect 39150 1492 39152 1532
rect 39152 1492 39194 1532
rect 39194 1492 39234 1532
rect 39234 1492 39274 1532
rect 39318 1492 39358 1532
rect 39358 1492 39398 1532
rect 39398 1492 39440 1532
rect 39440 1492 39442 1532
rect 39150 1450 39274 1492
rect 39318 1450 39442 1492
rect 51150 1532 51274 1574
rect 51318 1532 51442 1574
rect 51150 1492 51152 1532
rect 51152 1492 51194 1532
rect 51194 1492 51234 1532
rect 51234 1492 51274 1532
rect 51318 1492 51358 1532
rect 51358 1492 51398 1532
rect 51398 1492 51440 1532
rect 51440 1492 51442 1532
rect 51150 1450 51274 1492
rect 51318 1450 51442 1492
rect 63150 1532 63274 1574
rect 63318 1532 63442 1574
rect 63150 1492 63152 1532
rect 63152 1492 63194 1532
rect 63194 1492 63234 1532
rect 63234 1492 63274 1532
rect 63318 1492 63358 1532
rect 63358 1492 63398 1532
rect 63398 1492 63440 1532
rect 63440 1492 63442 1532
rect 63150 1450 63274 1492
rect 63318 1450 63442 1492
rect 75150 1532 75274 1574
rect 75318 1532 75442 1574
rect 75150 1492 75152 1532
rect 75152 1492 75194 1532
rect 75194 1492 75234 1532
rect 75234 1492 75274 1532
rect 75318 1492 75358 1532
rect 75358 1492 75398 1532
rect 75398 1492 75440 1532
rect 75440 1492 75442 1532
rect 75150 1450 75274 1492
rect 75318 1450 75442 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 16390 776 16514 818
rect 16558 776 16682 818
rect 16390 736 16392 776
rect 16392 736 16434 776
rect 16434 736 16474 776
rect 16474 736 16514 776
rect 16558 736 16598 776
rect 16598 736 16638 776
rect 16638 736 16680 776
rect 16680 736 16682 776
rect 16390 694 16514 736
rect 16558 694 16682 736
rect 28390 776 28514 818
rect 28558 776 28682 818
rect 28390 736 28392 776
rect 28392 736 28434 776
rect 28434 736 28474 776
rect 28474 736 28514 776
rect 28558 736 28598 776
rect 28598 736 28638 776
rect 28638 736 28680 776
rect 28680 736 28682 776
rect 28390 694 28514 736
rect 28558 694 28682 736
rect 40390 776 40514 818
rect 40558 776 40682 818
rect 40390 736 40392 776
rect 40392 736 40434 776
rect 40434 736 40474 776
rect 40474 736 40514 776
rect 40558 736 40598 776
rect 40598 736 40638 776
rect 40638 736 40680 776
rect 40680 736 40682 776
rect 40390 694 40514 736
rect 40558 694 40682 736
rect 52390 776 52514 818
rect 52558 776 52682 818
rect 52390 736 52392 776
rect 52392 736 52434 776
rect 52434 736 52474 776
rect 52474 736 52514 776
rect 52558 736 52598 776
rect 52598 736 52638 776
rect 52638 736 52680 776
rect 52680 736 52682 776
rect 52390 694 52514 736
rect 52558 694 52682 736
rect 64390 776 64514 818
rect 64558 776 64682 818
rect 64390 736 64392 776
rect 64392 736 64434 776
rect 64434 736 64474 776
rect 64474 736 64514 776
rect 64558 736 64598 776
rect 64598 736 64638 776
rect 64638 736 64680 776
rect 64680 736 64682 776
rect 64390 694 64514 736
rect 64558 694 64682 736
rect 76390 776 76514 818
rect 76558 776 76682 818
rect 76390 736 76392 776
rect 76392 736 76434 776
rect 76434 736 76474 776
rect 76474 736 76514 776
rect 76558 736 76598 776
rect 76598 736 76638 776
rect 76638 736 76680 776
rect 76680 736 76682 776
rect 76390 694 76514 736
rect 76558 694 76682 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 16316 38618 16756 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 15076 37862 15516 38600
rect 15076 37738 15150 37862
rect 15274 37738 15318 37862
rect 15442 37738 15516 37862
rect 15076 36350 15516 37738
rect 15076 36226 15150 36350
rect 15274 36226 15318 36350
rect 15442 36226 15516 36350
rect 15076 34838 15516 36226
rect 15076 34714 15150 34838
rect 15274 34714 15318 34838
rect 15442 34714 15516 34838
rect 15076 33326 15516 34714
rect 15076 33202 15150 33326
rect 15274 33202 15318 33326
rect 15442 33202 15516 33326
rect 15076 31814 15516 33202
rect 15076 31690 15150 31814
rect 15274 31690 15318 31814
rect 15442 31690 15516 31814
rect 15076 30302 15516 31690
rect 15076 30178 15150 30302
rect 15274 30178 15318 30302
rect 15442 30178 15516 30302
rect 15076 28790 15516 30178
rect 15076 28666 15150 28790
rect 15274 28666 15318 28790
rect 15442 28666 15516 28790
rect 15076 27278 15516 28666
rect 15076 27154 15150 27278
rect 15274 27154 15318 27278
rect 15442 27154 15516 27278
rect 15076 25766 15516 27154
rect 15076 25642 15150 25766
rect 15274 25642 15318 25766
rect 15442 25642 15516 25766
rect 15076 24254 15516 25642
rect 15076 24130 15150 24254
rect 15274 24130 15318 24254
rect 15442 24130 15516 24254
rect 15076 22742 15516 24130
rect 15076 22618 15150 22742
rect 15274 22618 15318 22742
rect 15442 22618 15516 22742
rect 15076 21230 15516 22618
rect 15076 21106 15150 21230
rect 15274 21106 15318 21230
rect 15442 21106 15516 21230
rect 15076 19718 15516 21106
rect 15076 19594 15150 19718
rect 15274 19594 15318 19718
rect 15442 19594 15516 19718
rect 15076 18206 15516 19594
rect 15076 18082 15150 18206
rect 15274 18082 15318 18206
rect 15442 18082 15516 18206
rect 15076 16694 15516 18082
rect 15076 16570 15150 16694
rect 15274 16570 15318 16694
rect 15442 16570 15516 16694
rect 15076 15182 15516 16570
rect 15076 15058 15150 15182
rect 15274 15058 15318 15182
rect 15442 15058 15516 15182
rect 15076 13670 15516 15058
rect 15076 13546 15150 13670
rect 15274 13546 15318 13670
rect 15442 13546 15516 13670
rect 15076 12158 15516 13546
rect 15076 12034 15150 12158
rect 15274 12034 15318 12158
rect 15442 12034 15516 12158
rect 15076 10646 15516 12034
rect 15076 10522 15150 10646
rect 15274 10522 15318 10646
rect 15442 10522 15516 10646
rect 15076 9134 15516 10522
rect 15076 9010 15150 9134
rect 15274 9010 15318 9134
rect 15442 9010 15516 9134
rect 15076 7622 15516 9010
rect 15076 7498 15150 7622
rect 15274 7498 15318 7622
rect 15442 7498 15516 7622
rect 15076 6110 15516 7498
rect 15076 5986 15150 6110
rect 15274 5986 15318 6110
rect 15442 5986 15516 6110
rect 15076 4598 15516 5986
rect 15076 4474 15150 4598
rect 15274 4474 15318 4598
rect 15442 4474 15516 4598
rect 15076 3086 15516 4474
rect 15076 2962 15150 3086
rect 15274 2962 15318 3086
rect 15442 2962 15516 3086
rect 15076 1574 15516 2962
rect 15076 1450 15150 1574
rect 15274 1450 15318 1574
rect 15442 1450 15516 1574
rect 15076 712 15516 1450
rect 16316 38494 16390 38618
rect 16514 38494 16558 38618
rect 16682 38494 16756 38618
rect 28316 38618 28756 38682
rect 16316 37106 16756 38494
rect 16316 36982 16390 37106
rect 16514 36982 16558 37106
rect 16682 36982 16756 37106
rect 16316 35594 16756 36982
rect 16316 35470 16390 35594
rect 16514 35470 16558 35594
rect 16682 35470 16756 35594
rect 16316 34082 16756 35470
rect 16316 33958 16390 34082
rect 16514 33958 16558 34082
rect 16682 33958 16756 34082
rect 16316 32570 16756 33958
rect 16316 32446 16390 32570
rect 16514 32446 16558 32570
rect 16682 32446 16756 32570
rect 16316 31058 16756 32446
rect 16316 30934 16390 31058
rect 16514 30934 16558 31058
rect 16682 30934 16756 31058
rect 16316 29546 16756 30934
rect 16316 29422 16390 29546
rect 16514 29422 16558 29546
rect 16682 29422 16756 29546
rect 16316 28034 16756 29422
rect 16316 27910 16390 28034
rect 16514 27910 16558 28034
rect 16682 27910 16756 28034
rect 16316 26522 16756 27910
rect 16316 26398 16390 26522
rect 16514 26398 16558 26522
rect 16682 26398 16756 26522
rect 16316 25010 16756 26398
rect 16316 24886 16390 25010
rect 16514 24886 16558 25010
rect 16682 24886 16756 25010
rect 16316 23498 16756 24886
rect 16316 23374 16390 23498
rect 16514 23374 16558 23498
rect 16682 23374 16756 23498
rect 16316 21986 16756 23374
rect 16316 21862 16390 21986
rect 16514 21862 16558 21986
rect 16682 21862 16756 21986
rect 16316 20474 16756 21862
rect 16316 20350 16390 20474
rect 16514 20350 16558 20474
rect 16682 20350 16756 20474
rect 16316 18962 16756 20350
rect 16316 18838 16390 18962
rect 16514 18838 16558 18962
rect 16682 18838 16756 18962
rect 16316 17450 16756 18838
rect 16316 17326 16390 17450
rect 16514 17326 16558 17450
rect 16682 17326 16756 17450
rect 16316 15938 16756 17326
rect 16316 15814 16390 15938
rect 16514 15814 16558 15938
rect 16682 15814 16756 15938
rect 16316 14426 16756 15814
rect 16316 14302 16390 14426
rect 16514 14302 16558 14426
rect 16682 14302 16756 14426
rect 16316 12914 16756 14302
rect 16316 12790 16390 12914
rect 16514 12790 16558 12914
rect 16682 12790 16756 12914
rect 16316 11402 16756 12790
rect 16316 11278 16390 11402
rect 16514 11278 16558 11402
rect 16682 11278 16756 11402
rect 16316 9890 16756 11278
rect 16316 9766 16390 9890
rect 16514 9766 16558 9890
rect 16682 9766 16756 9890
rect 16316 8378 16756 9766
rect 16316 8254 16390 8378
rect 16514 8254 16558 8378
rect 16682 8254 16756 8378
rect 16316 6866 16756 8254
rect 16316 6742 16390 6866
rect 16514 6742 16558 6866
rect 16682 6742 16756 6866
rect 16316 5354 16756 6742
rect 16316 5230 16390 5354
rect 16514 5230 16558 5354
rect 16682 5230 16756 5354
rect 16316 3842 16756 5230
rect 16316 3718 16390 3842
rect 16514 3718 16558 3842
rect 16682 3718 16756 3842
rect 16316 2330 16756 3718
rect 16316 2206 16390 2330
rect 16514 2206 16558 2330
rect 16682 2206 16756 2330
rect 16316 818 16756 2206
rect 4316 630 4756 694
rect 16316 694 16390 818
rect 16514 694 16558 818
rect 16682 694 16756 818
rect 27076 37862 27516 38600
rect 27076 37738 27150 37862
rect 27274 37738 27318 37862
rect 27442 37738 27516 37862
rect 27076 36350 27516 37738
rect 27076 36226 27150 36350
rect 27274 36226 27318 36350
rect 27442 36226 27516 36350
rect 27076 34838 27516 36226
rect 27076 34714 27150 34838
rect 27274 34714 27318 34838
rect 27442 34714 27516 34838
rect 27076 33326 27516 34714
rect 27076 33202 27150 33326
rect 27274 33202 27318 33326
rect 27442 33202 27516 33326
rect 27076 31814 27516 33202
rect 27076 31690 27150 31814
rect 27274 31690 27318 31814
rect 27442 31690 27516 31814
rect 27076 30302 27516 31690
rect 27076 30178 27150 30302
rect 27274 30178 27318 30302
rect 27442 30178 27516 30302
rect 27076 28790 27516 30178
rect 27076 28666 27150 28790
rect 27274 28666 27318 28790
rect 27442 28666 27516 28790
rect 27076 27278 27516 28666
rect 27076 27154 27150 27278
rect 27274 27154 27318 27278
rect 27442 27154 27516 27278
rect 27076 25766 27516 27154
rect 27076 25642 27150 25766
rect 27274 25642 27318 25766
rect 27442 25642 27516 25766
rect 27076 24254 27516 25642
rect 27076 24130 27150 24254
rect 27274 24130 27318 24254
rect 27442 24130 27516 24254
rect 27076 22742 27516 24130
rect 27076 22618 27150 22742
rect 27274 22618 27318 22742
rect 27442 22618 27516 22742
rect 27076 21230 27516 22618
rect 27076 21106 27150 21230
rect 27274 21106 27318 21230
rect 27442 21106 27516 21230
rect 27076 19718 27516 21106
rect 27076 19594 27150 19718
rect 27274 19594 27318 19718
rect 27442 19594 27516 19718
rect 27076 18206 27516 19594
rect 27076 18082 27150 18206
rect 27274 18082 27318 18206
rect 27442 18082 27516 18206
rect 27076 16694 27516 18082
rect 27076 16570 27150 16694
rect 27274 16570 27318 16694
rect 27442 16570 27516 16694
rect 27076 15182 27516 16570
rect 27076 15058 27150 15182
rect 27274 15058 27318 15182
rect 27442 15058 27516 15182
rect 27076 13670 27516 15058
rect 27076 13546 27150 13670
rect 27274 13546 27318 13670
rect 27442 13546 27516 13670
rect 27076 12158 27516 13546
rect 27076 12034 27150 12158
rect 27274 12034 27318 12158
rect 27442 12034 27516 12158
rect 27076 10646 27516 12034
rect 27076 10522 27150 10646
rect 27274 10522 27318 10646
rect 27442 10522 27516 10646
rect 27076 9134 27516 10522
rect 27076 9010 27150 9134
rect 27274 9010 27318 9134
rect 27442 9010 27516 9134
rect 27076 7622 27516 9010
rect 27076 7498 27150 7622
rect 27274 7498 27318 7622
rect 27442 7498 27516 7622
rect 27076 6110 27516 7498
rect 27076 5986 27150 6110
rect 27274 5986 27318 6110
rect 27442 5986 27516 6110
rect 27076 4598 27516 5986
rect 27076 4474 27150 4598
rect 27274 4474 27318 4598
rect 27442 4474 27516 4598
rect 27076 3086 27516 4474
rect 27076 2962 27150 3086
rect 27274 2962 27318 3086
rect 27442 2962 27516 3086
rect 27076 1574 27516 2962
rect 27076 1450 27150 1574
rect 27274 1450 27318 1574
rect 27442 1450 27516 1574
rect 27076 712 27516 1450
rect 28316 38494 28390 38618
rect 28514 38494 28558 38618
rect 28682 38494 28756 38618
rect 40316 38618 40756 38682
rect 28316 37106 28756 38494
rect 28316 36982 28390 37106
rect 28514 36982 28558 37106
rect 28682 36982 28756 37106
rect 28316 35594 28756 36982
rect 28316 35470 28390 35594
rect 28514 35470 28558 35594
rect 28682 35470 28756 35594
rect 28316 34082 28756 35470
rect 28316 33958 28390 34082
rect 28514 33958 28558 34082
rect 28682 33958 28756 34082
rect 28316 32570 28756 33958
rect 28316 32446 28390 32570
rect 28514 32446 28558 32570
rect 28682 32446 28756 32570
rect 28316 31058 28756 32446
rect 28316 30934 28390 31058
rect 28514 30934 28558 31058
rect 28682 30934 28756 31058
rect 28316 29546 28756 30934
rect 28316 29422 28390 29546
rect 28514 29422 28558 29546
rect 28682 29422 28756 29546
rect 28316 28034 28756 29422
rect 28316 27910 28390 28034
rect 28514 27910 28558 28034
rect 28682 27910 28756 28034
rect 28316 26522 28756 27910
rect 28316 26398 28390 26522
rect 28514 26398 28558 26522
rect 28682 26398 28756 26522
rect 28316 25010 28756 26398
rect 28316 24886 28390 25010
rect 28514 24886 28558 25010
rect 28682 24886 28756 25010
rect 28316 23498 28756 24886
rect 28316 23374 28390 23498
rect 28514 23374 28558 23498
rect 28682 23374 28756 23498
rect 28316 21986 28756 23374
rect 28316 21862 28390 21986
rect 28514 21862 28558 21986
rect 28682 21862 28756 21986
rect 28316 20474 28756 21862
rect 28316 20350 28390 20474
rect 28514 20350 28558 20474
rect 28682 20350 28756 20474
rect 28316 18962 28756 20350
rect 28316 18838 28390 18962
rect 28514 18838 28558 18962
rect 28682 18838 28756 18962
rect 28316 17450 28756 18838
rect 28316 17326 28390 17450
rect 28514 17326 28558 17450
rect 28682 17326 28756 17450
rect 28316 15938 28756 17326
rect 28316 15814 28390 15938
rect 28514 15814 28558 15938
rect 28682 15814 28756 15938
rect 28316 14426 28756 15814
rect 28316 14302 28390 14426
rect 28514 14302 28558 14426
rect 28682 14302 28756 14426
rect 28316 12914 28756 14302
rect 28316 12790 28390 12914
rect 28514 12790 28558 12914
rect 28682 12790 28756 12914
rect 28316 11402 28756 12790
rect 28316 11278 28390 11402
rect 28514 11278 28558 11402
rect 28682 11278 28756 11402
rect 28316 9890 28756 11278
rect 28316 9766 28390 9890
rect 28514 9766 28558 9890
rect 28682 9766 28756 9890
rect 28316 8378 28756 9766
rect 28316 8254 28390 8378
rect 28514 8254 28558 8378
rect 28682 8254 28756 8378
rect 28316 6866 28756 8254
rect 28316 6742 28390 6866
rect 28514 6742 28558 6866
rect 28682 6742 28756 6866
rect 28316 5354 28756 6742
rect 28316 5230 28390 5354
rect 28514 5230 28558 5354
rect 28682 5230 28756 5354
rect 28316 3842 28756 5230
rect 28316 3718 28390 3842
rect 28514 3718 28558 3842
rect 28682 3718 28756 3842
rect 28316 2330 28756 3718
rect 28316 2206 28390 2330
rect 28514 2206 28558 2330
rect 28682 2206 28756 2330
rect 28316 818 28756 2206
rect 16316 630 16756 694
rect 28316 694 28390 818
rect 28514 694 28558 818
rect 28682 694 28756 818
rect 39076 37862 39516 38600
rect 39076 37738 39150 37862
rect 39274 37738 39318 37862
rect 39442 37738 39516 37862
rect 39076 36350 39516 37738
rect 39076 36226 39150 36350
rect 39274 36226 39318 36350
rect 39442 36226 39516 36350
rect 39076 34838 39516 36226
rect 39076 34714 39150 34838
rect 39274 34714 39318 34838
rect 39442 34714 39516 34838
rect 39076 33326 39516 34714
rect 39076 33202 39150 33326
rect 39274 33202 39318 33326
rect 39442 33202 39516 33326
rect 39076 31814 39516 33202
rect 39076 31690 39150 31814
rect 39274 31690 39318 31814
rect 39442 31690 39516 31814
rect 39076 30302 39516 31690
rect 39076 30178 39150 30302
rect 39274 30178 39318 30302
rect 39442 30178 39516 30302
rect 39076 28790 39516 30178
rect 39076 28666 39150 28790
rect 39274 28666 39318 28790
rect 39442 28666 39516 28790
rect 39076 27278 39516 28666
rect 39076 27154 39150 27278
rect 39274 27154 39318 27278
rect 39442 27154 39516 27278
rect 39076 25766 39516 27154
rect 39076 25642 39150 25766
rect 39274 25642 39318 25766
rect 39442 25642 39516 25766
rect 39076 24254 39516 25642
rect 39076 24130 39150 24254
rect 39274 24130 39318 24254
rect 39442 24130 39516 24254
rect 39076 22742 39516 24130
rect 39076 22618 39150 22742
rect 39274 22618 39318 22742
rect 39442 22618 39516 22742
rect 39076 21230 39516 22618
rect 39076 21106 39150 21230
rect 39274 21106 39318 21230
rect 39442 21106 39516 21230
rect 39076 19718 39516 21106
rect 39076 19594 39150 19718
rect 39274 19594 39318 19718
rect 39442 19594 39516 19718
rect 39076 18206 39516 19594
rect 39076 18082 39150 18206
rect 39274 18082 39318 18206
rect 39442 18082 39516 18206
rect 39076 16694 39516 18082
rect 39076 16570 39150 16694
rect 39274 16570 39318 16694
rect 39442 16570 39516 16694
rect 39076 15182 39516 16570
rect 39076 15058 39150 15182
rect 39274 15058 39318 15182
rect 39442 15058 39516 15182
rect 39076 13670 39516 15058
rect 39076 13546 39150 13670
rect 39274 13546 39318 13670
rect 39442 13546 39516 13670
rect 39076 12158 39516 13546
rect 39076 12034 39150 12158
rect 39274 12034 39318 12158
rect 39442 12034 39516 12158
rect 39076 10646 39516 12034
rect 39076 10522 39150 10646
rect 39274 10522 39318 10646
rect 39442 10522 39516 10646
rect 39076 9134 39516 10522
rect 39076 9010 39150 9134
rect 39274 9010 39318 9134
rect 39442 9010 39516 9134
rect 39076 7622 39516 9010
rect 39076 7498 39150 7622
rect 39274 7498 39318 7622
rect 39442 7498 39516 7622
rect 39076 6110 39516 7498
rect 39076 5986 39150 6110
rect 39274 5986 39318 6110
rect 39442 5986 39516 6110
rect 39076 4598 39516 5986
rect 39076 4474 39150 4598
rect 39274 4474 39318 4598
rect 39442 4474 39516 4598
rect 39076 3086 39516 4474
rect 39076 2962 39150 3086
rect 39274 2962 39318 3086
rect 39442 2962 39516 3086
rect 39076 1574 39516 2962
rect 39076 1450 39150 1574
rect 39274 1450 39318 1574
rect 39442 1450 39516 1574
rect 39076 712 39516 1450
rect 40316 38494 40390 38618
rect 40514 38494 40558 38618
rect 40682 38494 40756 38618
rect 52316 38618 52756 38682
rect 40316 37106 40756 38494
rect 40316 36982 40390 37106
rect 40514 36982 40558 37106
rect 40682 36982 40756 37106
rect 40316 35594 40756 36982
rect 40316 35470 40390 35594
rect 40514 35470 40558 35594
rect 40682 35470 40756 35594
rect 40316 34082 40756 35470
rect 40316 33958 40390 34082
rect 40514 33958 40558 34082
rect 40682 33958 40756 34082
rect 40316 32570 40756 33958
rect 40316 32446 40390 32570
rect 40514 32446 40558 32570
rect 40682 32446 40756 32570
rect 40316 31058 40756 32446
rect 40316 30934 40390 31058
rect 40514 30934 40558 31058
rect 40682 30934 40756 31058
rect 40316 29546 40756 30934
rect 40316 29422 40390 29546
rect 40514 29422 40558 29546
rect 40682 29422 40756 29546
rect 40316 28034 40756 29422
rect 40316 27910 40390 28034
rect 40514 27910 40558 28034
rect 40682 27910 40756 28034
rect 40316 26522 40756 27910
rect 40316 26398 40390 26522
rect 40514 26398 40558 26522
rect 40682 26398 40756 26522
rect 40316 25010 40756 26398
rect 40316 24886 40390 25010
rect 40514 24886 40558 25010
rect 40682 24886 40756 25010
rect 40316 23498 40756 24886
rect 40316 23374 40390 23498
rect 40514 23374 40558 23498
rect 40682 23374 40756 23498
rect 40316 21986 40756 23374
rect 40316 21862 40390 21986
rect 40514 21862 40558 21986
rect 40682 21862 40756 21986
rect 40316 20474 40756 21862
rect 40316 20350 40390 20474
rect 40514 20350 40558 20474
rect 40682 20350 40756 20474
rect 40316 18962 40756 20350
rect 40316 18838 40390 18962
rect 40514 18838 40558 18962
rect 40682 18838 40756 18962
rect 40316 17450 40756 18838
rect 40316 17326 40390 17450
rect 40514 17326 40558 17450
rect 40682 17326 40756 17450
rect 40316 15938 40756 17326
rect 40316 15814 40390 15938
rect 40514 15814 40558 15938
rect 40682 15814 40756 15938
rect 40316 14426 40756 15814
rect 40316 14302 40390 14426
rect 40514 14302 40558 14426
rect 40682 14302 40756 14426
rect 40316 12914 40756 14302
rect 40316 12790 40390 12914
rect 40514 12790 40558 12914
rect 40682 12790 40756 12914
rect 40316 11402 40756 12790
rect 40316 11278 40390 11402
rect 40514 11278 40558 11402
rect 40682 11278 40756 11402
rect 40316 9890 40756 11278
rect 40316 9766 40390 9890
rect 40514 9766 40558 9890
rect 40682 9766 40756 9890
rect 40316 8378 40756 9766
rect 40316 8254 40390 8378
rect 40514 8254 40558 8378
rect 40682 8254 40756 8378
rect 40316 6866 40756 8254
rect 40316 6742 40390 6866
rect 40514 6742 40558 6866
rect 40682 6742 40756 6866
rect 40316 5354 40756 6742
rect 40316 5230 40390 5354
rect 40514 5230 40558 5354
rect 40682 5230 40756 5354
rect 40316 3842 40756 5230
rect 40316 3718 40390 3842
rect 40514 3718 40558 3842
rect 40682 3718 40756 3842
rect 40316 2330 40756 3718
rect 40316 2206 40390 2330
rect 40514 2206 40558 2330
rect 40682 2206 40756 2330
rect 40316 818 40756 2206
rect 28316 630 28756 694
rect 40316 694 40390 818
rect 40514 694 40558 818
rect 40682 694 40756 818
rect 51076 37862 51516 38600
rect 51076 37738 51150 37862
rect 51274 37738 51318 37862
rect 51442 37738 51516 37862
rect 51076 36350 51516 37738
rect 51076 36226 51150 36350
rect 51274 36226 51318 36350
rect 51442 36226 51516 36350
rect 51076 34838 51516 36226
rect 51076 34714 51150 34838
rect 51274 34714 51318 34838
rect 51442 34714 51516 34838
rect 51076 33326 51516 34714
rect 51076 33202 51150 33326
rect 51274 33202 51318 33326
rect 51442 33202 51516 33326
rect 51076 31814 51516 33202
rect 51076 31690 51150 31814
rect 51274 31690 51318 31814
rect 51442 31690 51516 31814
rect 51076 30302 51516 31690
rect 51076 30178 51150 30302
rect 51274 30178 51318 30302
rect 51442 30178 51516 30302
rect 51076 28790 51516 30178
rect 51076 28666 51150 28790
rect 51274 28666 51318 28790
rect 51442 28666 51516 28790
rect 51076 27278 51516 28666
rect 51076 27154 51150 27278
rect 51274 27154 51318 27278
rect 51442 27154 51516 27278
rect 51076 25766 51516 27154
rect 51076 25642 51150 25766
rect 51274 25642 51318 25766
rect 51442 25642 51516 25766
rect 51076 15182 51516 25642
rect 51076 15058 51150 15182
rect 51274 15058 51318 15182
rect 51442 15058 51516 15182
rect 51076 13670 51516 15058
rect 51076 13546 51150 13670
rect 51274 13546 51318 13670
rect 51442 13546 51516 13670
rect 51076 12158 51516 13546
rect 51076 12034 51150 12158
rect 51274 12034 51318 12158
rect 51442 12034 51516 12158
rect 51076 10646 51516 12034
rect 51076 10522 51150 10646
rect 51274 10522 51318 10646
rect 51442 10522 51516 10646
rect 51076 9134 51516 10522
rect 51076 9010 51150 9134
rect 51274 9010 51318 9134
rect 51442 9010 51516 9134
rect 51076 7622 51516 9010
rect 51076 7498 51150 7622
rect 51274 7498 51318 7622
rect 51442 7498 51516 7622
rect 51076 6110 51516 7498
rect 51076 5986 51150 6110
rect 51274 5986 51318 6110
rect 51442 5986 51516 6110
rect 51076 4598 51516 5986
rect 51076 4474 51150 4598
rect 51274 4474 51318 4598
rect 51442 4474 51516 4598
rect 51076 3086 51516 4474
rect 51076 2962 51150 3086
rect 51274 2962 51318 3086
rect 51442 2962 51516 3086
rect 51076 1574 51516 2962
rect 51076 1450 51150 1574
rect 51274 1450 51318 1574
rect 51442 1450 51516 1574
rect 51076 712 51516 1450
rect 52316 38494 52390 38618
rect 52514 38494 52558 38618
rect 52682 38494 52756 38618
rect 64316 38618 64756 38682
rect 52316 37106 52756 38494
rect 52316 36982 52390 37106
rect 52514 36982 52558 37106
rect 52682 36982 52756 37106
rect 52316 35594 52756 36982
rect 52316 35470 52390 35594
rect 52514 35470 52558 35594
rect 52682 35470 52756 35594
rect 52316 34082 52756 35470
rect 52316 33958 52390 34082
rect 52514 33958 52558 34082
rect 52682 33958 52756 34082
rect 52316 32570 52756 33958
rect 52316 32446 52390 32570
rect 52514 32446 52558 32570
rect 52682 32446 52756 32570
rect 52316 31058 52756 32446
rect 52316 30934 52390 31058
rect 52514 30934 52558 31058
rect 52682 30934 52756 31058
rect 52316 29546 52756 30934
rect 52316 29422 52390 29546
rect 52514 29422 52558 29546
rect 52682 29422 52756 29546
rect 52316 28034 52756 29422
rect 52316 27910 52390 28034
rect 52514 27910 52558 28034
rect 52682 27910 52756 28034
rect 52316 26522 52756 27910
rect 52316 26398 52390 26522
rect 52514 26398 52558 26522
rect 52682 26398 52756 26522
rect 52316 25010 52756 26398
rect 52316 24886 52390 25010
rect 52514 24886 52558 25010
rect 52682 24886 52756 25010
rect 52316 14426 52756 24886
rect 52316 14302 52390 14426
rect 52514 14302 52558 14426
rect 52682 14302 52756 14426
rect 52316 12914 52756 14302
rect 52316 12790 52390 12914
rect 52514 12790 52558 12914
rect 52682 12790 52756 12914
rect 52316 11402 52756 12790
rect 52316 11278 52390 11402
rect 52514 11278 52558 11402
rect 52682 11278 52756 11402
rect 52316 9890 52756 11278
rect 52316 9766 52390 9890
rect 52514 9766 52558 9890
rect 52682 9766 52756 9890
rect 52316 8378 52756 9766
rect 52316 8254 52390 8378
rect 52514 8254 52558 8378
rect 52682 8254 52756 8378
rect 52316 6866 52756 8254
rect 52316 6742 52390 6866
rect 52514 6742 52558 6866
rect 52682 6742 52756 6866
rect 52316 5354 52756 6742
rect 52316 5230 52390 5354
rect 52514 5230 52558 5354
rect 52682 5230 52756 5354
rect 52316 3842 52756 5230
rect 52316 3718 52390 3842
rect 52514 3718 52558 3842
rect 52682 3718 52756 3842
rect 52316 2330 52756 3718
rect 52316 2206 52390 2330
rect 52514 2206 52558 2330
rect 52682 2206 52756 2330
rect 52316 818 52756 2206
rect 40316 630 40756 694
rect 52316 694 52390 818
rect 52514 694 52558 818
rect 52682 694 52756 818
rect 63076 37862 63516 38600
rect 63076 37738 63150 37862
rect 63274 37738 63318 37862
rect 63442 37738 63516 37862
rect 63076 36350 63516 37738
rect 63076 36226 63150 36350
rect 63274 36226 63318 36350
rect 63442 36226 63516 36350
rect 63076 34838 63516 36226
rect 63076 34714 63150 34838
rect 63274 34714 63318 34838
rect 63442 34714 63516 34838
rect 63076 33326 63516 34714
rect 63076 33202 63150 33326
rect 63274 33202 63318 33326
rect 63442 33202 63516 33326
rect 63076 31814 63516 33202
rect 63076 31690 63150 31814
rect 63274 31690 63318 31814
rect 63442 31690 63516 31814
rect 63076 30302 63516 31690
rect 63076 30178 63150 30302
rect 63274 30178 63318 30302
rect 63442 30178 63516 30302
rect 63076 28790 63516 30178
rect 63076 28666 63150 28790
rect 63274 28666 63318 28790
rect 63442 28666 63516 28790
rect 63076 27278 63516 28666
rect 63076 27154 63150 27278
rect 63274 27154 63318 27278
rect 63442 27154 63516 27278
rect 63076 25766 63516 27154
rect 63076 25642 63150 25766
rect 63274 25642 63318 25766
rect 63442 25642 63516 25766
rect 63076 19665 63516 25642
rect 63076 19541 63150 19665
rect 63274 19541 63318 19665
rect 63442 19541 63516 19665
rect 63076 19497 63516 19541
rect 63076 19373 63150 19497
rect 63274 19373 63318 19497
rect 63442 19373 63516 19497
rect 63076 19329 63516 19373
rect 63076 19205 63150 19329
rect 63274 19205 63318 19329
rect 63442 19205 63516 19329
rect 63076 19161 63516 19205
rect 63076 19037 63150 19161
rect 63274 19037 63318 19161
rect 63442 19037 63516 19161
rect 63076 18993 63516 19037
rect 63076 18869 63150 18993
rect 63274 18869 63318 18993
rect 63442 18869 63516 18993
rect 63076 18825 63516 18869
rect 63076 18701 63150 18825
rect 63274 18701 63318 18825
rect 63442 18701 63516 18825
rect 63076 18657 63516 18701
rect 63076 18533 63150 18657
rect 63274 18533 63318 18657
rect 63442 18533 63516 18657
rect 63076 18489 63516 18533
rect 63076 18365 63150 18489
rect 63274 18365 63318 18489
rect 63442 18365 63516 18489
rect 63076 18321 63516 18365
rect 63076 18197 63150 18321
rect 63274 18197 63318 18321
rect 63442 18197 63516 18321
rect 63076 18153 63516 18197
rect 63076 18029 63150 18153
rect 63274 18029 63318 18153
rect 63442 18029 63516 18153
rect 63076 17985 63516 18029
rect 63076 17861 63150 17985
rect 63274 17861 63318 17985
rect 63442 17861 63516 17985
rect 63076 17817 63516 17861
rect 63076 17693 63150 17817
rect 63274 17693 63318 17817
rect 63442 17693 63516 17817
rect 63076 17649 63516 17693
rect 63076 17525 63150 17649
rect 63274 17525 63318 17649
rect 63442 17525 63516 17649
rect 63076 15182 63516 17525
rect 63076 15058 63150 15182
rect 63274 15058 63318 15182
rect 63442 15058 63516 15182
rect 63076 13670 63516 15058
rect 63076 13546 63150 13670
rect 63274 13546 63318 13670
rect 63442 13546 63516 13670
rect 63076 12158 63516 13546
rect 63076 12034 63150 12158
rect 63274 12034 63318 12158
rect 63442 12034 63516 12158
rect 63076 10646 63516 12034
rect 63076 10522 63150 10646
rect 63274 10522 63318 10646
rect 63442 10522 63516 10646
rect 63076 9134 63516 10522
rect 63076 9010 63150 9134
rect 63274 9010 63318 9134
rect 63442 9010 63516 9134
rect 63076 7622 63516 9010
rect 63076 7498 63150 7622
rect 63274 7498 63318 7622
rect 63442 7498 63516 7622
rect 63076 6110 63516 7498
rect 63076 5986 63150 6110
rect 63274 5986 63318 6110
rect 63442 5986 63516 6110
rect 63076 4598 63516 5986
rect 63076 4474 63150 4598
rect 63274 4474 63318 4598
rect 63442 4474 63516 4598
rect 63076 3086 63516 4474
rect 63076 2962 63150 3086
rect 63274 2962 63318 3086
rect 63442 2962 63516 3086
rect 63076 1574 63516 2962
rect 63076 1450 63150 1574
rect 63274 1450 63318 1574
rect 63442 1450 63516 1574
rect 63076 712 63516 1450
rect 64316 38494 64390 38618
rect 64514 38494 64558 38618
rect 64682 38494 64756 38618
rect 76316 38618 76756 38682
rect 64316 37106 64756 38494
rect 64316 36982 64390 37106
rect 64514 36982 64558 37106
rect 64682 36982 64756 37106
rect 64316 35594 64756 36982
rect 64316 35470 64390 35594
rect 64514 35470 64558 35594
rect 64682 35470 64756 35594
rect 64316 34082 64756 35470
rect 64316 33958 64390 34082
rect 64514 33958 64558 34082
rect 64682 33958 64756 34082
rect 64316 32570 64756 33958
rect 64316 32446 64390 32570
rect 64514 32446 64558 32570
rect 64682 32446 64756 32570
rect 64316 31058 64756 32446
rect 64316 30934 64390 31058
rect 64514 30934 64558 31058
rect 64682 30934 64756 31058
rect 64316 29546 64756 30934
rect 64316 29422 64390 29546
rect 64514 29422 64558 29546
rect 64682 29422 64756 29546
rect 64316 28034 64756 29422
rect 64316 27910 64390 28034
rect 64514 27910 64558 28034
rect 64682 27910 64756 28034
rect 64316 26522 64756 27910
rect 64316 26398 64390 26522
rect 64514 26398 64558 26522
rect 64682 26398 64756 26522
rect 64316 25010 64756 26398
rect 64316 24886 64390 25010
rect 64514 24886 64558 25010
rect 64682 24886 64756 25010
rect 64316 22541 64756 24886
rect 64316 22417 64390 22541
rect 64514 22417 64558 22541
rect 64682 22417 64756 22541
rect 64316 22373 64756 22417
rect 64316 22249 64390 22373
rect 64514 22249 64558 22373
rect 64682 22249 64756 22373
rect 64316 22205 64756 22249
rect 64316 22081 64390 22205
rect 64514 22081 64558 22205
rect 64682 22081 64756 22205
rect 64316 22037 64756 22081
rect 64316 21913 64390 22037
rect 64514 21913 64558 22037
rect 64682 21913 64756 22037
rect 64316 21869 64756 21913
rect 64316 21745 64390 21869
rect 64514 21745 64558 21869
rect 64682 21745 64756 21869
rect 64316 21701 64756 21745
rect 64316 21577 64390 21701
rect 64514 21577 64558 21701
rect 64682 21577 64756 21701
rect 64316 21533 64756 21577
rect 64316 21409 64390 21533
rect 64514 21409 64558 21533
rect 64682 21409 64756 21533
rect 64316 21365 64756 21409
rect 64316 21241 64390 21365
rect 64514 21241 64558 21365
rect 64682 21241 64756 21365
rect 64316 21197 64756 21241
rect 64316 21073 64390 21197
rect 64514 21073 64558 21197
rect 64682 21073 64756 21197
rect 64316 21029 64756 21073
rect 64316 20905 64390 21029
rect 64514 20905 64558 21029
rect 64682 20905 64756 21029
rect 64316 20861 64756 20905
rect 64316 20737 64390 20861
rect 64514 20737 64558 20861
rect 64682 20737 64756 20861
rect 64316 20693 64756 20737
rect 64316 20569 64390 20693
rect 64514 20569 64558 20693
rect 64682 20569 64756 20693
rect 64316 20525 64756 20569
rect 64316 20401 64390 20525
rect 64514 20401 64558 20525
rect 64682 20401 64756 20525
rect 64316 14426 64756 20401
rect 64316 14302 64390 14426
rect 64514 14302 64558 14426
rect 64682 14302 64756 14426
rect 64316 12914 64756 14302
rect 64316 12790 64390 12914
rect 64514 12790 64558 12914
rect 64682 12790 64756 12914
rect 64316 11402 64756 12790
rect 64316 11278 64390 11402
rect 64514 11278 64558 11402
rect 64682 11278 64756 11402
rect 64316 9890 64756 11278
rect 64316 9766 64390 9890
rect 64514 9766 64558 9890
rect 64682 9766 64756 9890
rect 64316 8378 64756 9766
rect 64316 8254 64390 8378
rect 64514 8254 64558 8378
rect 64682 8254 64756 8378
rect 64316 6866 64756 8254
rect 64316 6742 64390 6866
rect 64514 6742 64558 6866
rect 64682 6742 64756 6866
rect 64316 5354 64756 6742
rect 64316 5230 64390 5354
rect 64514 5230 64558 5354
rect 64682 5230 64756 5354
rect 64316 3842 64756 5230
rect 64316 3718 64390 3842
rect 64514 3718 64558 3842
rect 64682 3718 64756 3842
rect 64316 2330 64756 3718
rect 64316 2206 64390 2330
rect 64514 2206 64558 2330
rect 64682 2206 64756 2330
rect 64316 818 64756 2206
rect 52316 630 52756 694
rect 64316 694 64390 818
rect 64514 694 64558 818
rect 64682 694 64756 818
rect 75076 37862 75516 38600
rect 75076 37738 75150 37862
rect 75274 37738 75318 37862
rect 75442 37738 75516 37862
rect 75076 36350 75516 37738
rect 75076 36226 75150 36350
rect 75274 36226 75318 36350
rect 75442 36226 75516 36350
rect 75076 34838 75516 36226
rect 75076 34714 75150 34838
rect 75274 34714 75318 34838
rect 75442 34714 75516 34838
rect 75076 33326 75516 34714
rect 75076 33202 75150 33326
rect 75274 33202 75318 33326
rect 75442 33202 75516 33326
rect 75076 31814 75516 33202
rect 75076 31690 75150 31814
rect 75274 31690 75318 31814
rect 75442 31690 75516 31814
rect 75076 30302 75516 31690
rect 75076 30178 75150 30302
rect 75274 30178 75318 30302
rect 75442 30178 75516 30302
rect 75076 28790 75516 30178
rect 75076 28666 75150 28790
rect 75274 28666 75318 28790
rect 75442 28666 75516 28790
rect 75076 27278 75516 28666
rect 75076 27154 75150 27278
rect 75274 27154 75318 27278
rect 75442 27154 75516 27278
rect 75076 25766 75516 27154
rect 75076 25642 75150 25766
rect 75274 25642 75318 25766
rect 75442 25642 75516 25766
rect 75076 19665 75516 25642
rect 75076 19541 75150 19665
rect 75274 19541 75318 19665
rect 75442 19541 75516 19665
rect 75076 19497 75516 19541
rect 75076 19373 75150 19497
rect 75274 19373 75318 19497
rect 75442 19373 75516 19497
rect 75076 19329 75516 19373
rect 75076 19205 75150 19329
rect 75274 19205 75318 19329
rect 75442 19205 75516 19329
rect 75076 19161 75516 19205
rect 75076 19037 75150 19161
rect 75274 19037 75318 19161
rect 75442 19037 75516 19161
rect 75076 18993 75516 19037
rect 75076 18869 75150 18993
rect 75274 18869 75318 18993
rect 75442 18869 75516 18993
rect 75076 18825 75516 18869
rect 75076 18701 75150 18825
rect 75274 18701 75318 18825
rect 75442 18701 75516 18825
rect 75076 18657 75516 18701
rect 75076 18533 75150 18657
rect 75274 18533 75318 18657
rect 75442 18533 75516 18657
rect 75076 18489 75516 18533
rect 75076 18365 75150 18489
rect 75274 18365 75318 18489
rect 75442 18365 75516 18489
rect 75076 18321 75516 18365
rect 75076 18197 75150 18321
rect 75274 18197 75318 18321
rect 75442 18197 75516 18321
rect 75076 18153 75516 18197
rect 75076 18029 75150 18153
rect 75274 18029 75318 18153
rect 75442 18029 75516 18153
rect 75076 17985 75516 18029
rect 75076 17861 75150 17985
rect 75274 17861 75318 17985
rect 75442 17861 75516 17985
rect 75076 17817 75516 17861
rect 75076 17693 75150 17817
rect 75274 17693 75318 17817
rect 75442 17693 75516 17817
rect 75076 17649 75516 17693
rect 75076 17525 75150 17649
rect 75274 17525 75318 17649
rect 75442 17525 75516 17649
rect 75076 15182 75516 17525
rect 75076 15058 75150 15182
rect 75274 15058 75318 15182
rect 75442 15058 75516 15182
rect 75076 13670 75516 15058
rect 75076 13546 75150 13670
rect 75274 13546 75318 13670
rect 75442 13546 75516 13670
rect 75076 12158 75516 13546
rect 75076 12034 75150 12158
rect 75274 12034 75318 12158
rect 75442 12034 75516 12158
rect 75076 10646 75516 12034
rect 75076 10522 75150 10646
rect 75274 10522 75318 10646
rect 75442 10522 75516 10646
rect 75076 9134 75516 10522
rect 75076 9010 75150 9134
rect 75274 9010 75318 9134
rect 75442 9010 75516 9134
rect 75076 7622 75516 9010
rect 75076 7498 75150 7622
rect 75274 7498 75318 7622
rect 75442 7498 75516 7622
rect 75076 6110 75516 7498
rect 75076 5986 75150 6110
rect 75274 5986 75318 6110
rect 75442 5986 75516 6110
rect 75076 4598 75516 5986
rect 75076 4474 75150 4598
rect 75274 4474 75318 4598
rect 75442 4474 75516 4598
rect 75076 3086 75516 4474
rect 75076 2962 75150 3086
rect 75274 2962 75318 3086
rect 75442 2962 75516 3086
rect 75076 1574 75516 2962
rect 75076 1450 75150 1574
rect 75274 1450 75318 1574
rect 75442 1450 75516 1574
rect 75076 712 75516 1450
rect 76316 38494 76390 38618
rect 76514 38494 76558 38618
rect 76682 38494 76756 38618
rect 76316 37106 76756 38494
rect 76316 36982 76390 37106
rect 76514 36982 76558 37106
rect 76682 36982 76756 37106
rect 76316 35594 76756 36982
rect 76316 35470 76390 35594
rect 76514 35470 76558 35594
rect 76682 35470 76756 35594
rect 76316 34082 76756 35470
rect 76316 33958 76390 34082
rect 76514 33958 76558 34082
rect 76682 33958 76756 34082
rect 76316 32570 76756 33958
rect 76316 32446 76390 32570
rect 76514 32446 76558 32570
rect 76682 32446 76756 32570
rect 76316 31058 76756 32446
rect 76316 30934 76390 31058
rect 76514 30934 76558 31058
rect 76682 30934 76756 31058
rect 76316 29546 76756 30934
rect 76316 29422 76390 29546
rect 76514 29422 76558 29546
rect 76682 29422 76756 29546
rect 76316 28034 76756 29422
rect 76316 27910 76390 28034
rect 76514 27910 76558 28034
rect 76682 27910 76756 28034
rect 76316 26522 76756 27910
rect 76316 26398 76390 26522
rect 76514 26398 76558 26522
rect 76682 26398 76756 26522
rect 76316 25010 76756 26398
rect 76316 24886 76390 25010
rect 76514 24886 76558 25010
rect 76682 24886 76756 25010
rect 76316 22541 76756 24886
rect 76316 22417 76390 22541
rect 76514 22417 76558 22541
rect 76682 22417 76756 22541
rect 76316 22373 76756 22417
rect 76316 22249 76390 22373
rect 76514 22249 76558 22373
rect 76682 22249 76756 22373
rect 76316 22205 76756 22249
rect 76316 22081 76390 22205
rect 76514 22081 76558 22205
rect 76682 22081 76756 22205
rect 76316 22037 76756 22081
rect 76316 21913 76390 22037
rect 76514 21913 76558 22037
rect 76682 21913 76756 22037
rect 76316 21869 76756 21913
rect 76316 21745 76390 21869
rect 76514 21745 76558 21869
rect 76682 21745 76756 21869
rect 76316 21701 76756 21745
rect 76316 21577 76390 21701
rect 76514 21577 76558 21701
rect 76682 21577 76756 21701
rect 76316 21533 76756 21577
rect 76316 21409 76390 21533
rect 76514 21409 76558 21533
rect 76682 21409 76756 21533
rect 76316 21365 76756 21409
rect 76316 21241 76390 21365
rect 76514 21241 76558 21365
rect 76682 21241 76756 21365
rect 76316 21197 76756 21241
rect 76316 21073 76390 21197
rect 76514 21073 76558 21197
rect 76682 21073 76756 21197
rect 76316 21029 76756 21073
rect 76316 20905 76390 21029
rect 76514 20905 76558 21029
rect 76682 20905 76756 21029
rect 76316 20861 76756 20905
rect 76316 20737 76390 20861
rect 76514 20737 76558 20861
rect 76682 20737 76756 20861
rect 76316 20693 76756 20737
rect 76316 20569 76390 20693
rect 76514 20569 76558 20693
rect 76682 20569 76756 20693
rect 76316 20525 76756 20569
rect 76316 20401 76390 20525
rect 76514 20401 76558 20525
rect 76682 20401 76756 20525
rect 76316 14426 76756 20401
rect 78596 23834 78924 23936
rect 78596 23710 78698 23834
rect 78822 23710 78924 23834
rect 78596 16274 78924 23710
rect 78596 16150 78698 16274
rect 78822 16150 78924 16274
rect 78596 16048 78924 16150
rect 76316 14302 76390 14426
rect 76514 14302 76558 14426
rect 76682 14302 76756 14426
rect 76316 12914 76756 14302
rect 76316 12790 76390 12914
rect 76514 12790 76558 12914
rect 76682 12790 76756 12914
rect 76316 11402 76756 12790
rect 76316 11278 76390 11402
rect 76514 11278 76558 11402
rect 76682 11278 76756 11402
rect 76316 9890 76756 11278
rect 76316 9766 76390 9890
rect 76514 9766 76558 9890
rect 76682 9766 76756 9890
rect 76316 8378 76756 9766
rect 76316 8254 76390 8378
rect 76514 8254 76558 8378
rect 76682 8254 76756 8378
rect 76316 6866 76756 8254
rect 76316 6742 76390 6866
rect 76514 6742 76558 6866
rect 76682 6742 76756 6866
rect 76316 5354 76756 6742
rect 76316 5230 76390 5354
rect 76514 5230 76558 5354
rect 76682 5230 76756 5354
rect 76316 3842 76756 5230
rect 76316 3718 76390 3842
rect 76514 3718 76558 3842
rect 76682 3718 76756 3842
rect 76316 2330 76756 3718
rect 76316 2206 76390 2330
rect 76514 2206 76558 2330
rect 76682 2206 76756 2330
rect 76316 818 76756 2206
rect 64316 630 64756 694
rect 76316 694 76390 818
rect 76514 694 76558 818
rect 76682 694 76756 818
rect 76316 630 76756 694
use sg13g2_inv_1  _1284_
timestamp 1676382929
transform 1 0 52224 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1285_
timestamp 1676382929
transform 1 0 3648 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1286_
timestamp 1676382929
transform 1 0 52512 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1287_
timestamp 1676382929
transform 1 0 52512 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1288_
timestamp 1676382929
transform 1 0 54720 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1289_
timestamp 1676382929
transform 1 0 55008 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1290_
timestamp 1676382929
transform 1 0 55776 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1291_
timestamp 1676382929
transform 1 0 56064 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1292_
timestamp 1676382929
transform 1 0 56352 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1293_
timestamp 1676382929
transform 1 0 56736 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1294_
timestamp 1676382929
transform 1 0 57216 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1295_
timestamp 1676382929
transform 1 0 57600 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1296_
timestamp 1676382929
transform 1 0 57984 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1297_
timestamp 1676382929
transform 1 0 58368 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1298_
timestamp 1676382929
transform 1 0 58848 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1299_
timestamp 1676382929
transform 1 0 59232 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1300_
timestamp 1676382929
transform 1 0 59616 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1301_
timestamp 1676382929
transform 1 0 60000 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1302_
timestamp 1676382929
transform 1 0 60384 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1303_
timestamp 1676382929
transform 1 0 60768 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1304_
timestamp 1676382929
transform 1 0 61248 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1305_
timestamp 1676382929
transform 1 0 61632 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1306_
timestamp 1676382929
transform 1 0 62016 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1307_
timestamp 1676382929
transform 1 0 62400 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1308_
timestamp 1676382929
transform 1 0 62784 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1309_
timestamp 1676382929
transform 1 0 63168 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1310_
timestamp 1676382929
transform 1 0 63648 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1311_
timestamp 1676382929
transform 1 0 64032 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1312_
timestamp 1676382929
transform 1 0 64416 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1313_
timestamp 1676382929
transform 1 0 64800 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1314_
timestamp 1676382929
transform 1 0 65184 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1315_
timestamp 1676382929
transform 1 0 65664 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1316_
timestamp 1676382929
transform 1 0 66048 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1317_
timestamp 1676382929
transform 1 0 66432 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1318_
timestamp 1676382929
transform 1 0 66816 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1319_
timestamp 1676382929
transform 1 0 67200 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1320_
timestamp 1676382929
transform 1 0 67680 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1321_
timestamp 1676382929
transform 1 0 68064 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1322_
timestamp 1676382929
transform 1 0 68448 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1323_
timestamp 1676382929
transform 1 0 68832 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1324_
timestamp 1676382929
transform 1 0 69216 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1325_
timestamp 1676382929
transform 1 0 69696 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1326_
timestamp 1676382929
transform 1 0 70080 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1327_
timestamp 1676382929
transform 1 0 70464 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1328_
timestamp 1676382929
transform 1 0 70848 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1329_
timestamp 1676382929
transform 1 0 71232 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1330_
timestamp 1676382929
transform 1 0 71616 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1331_
timestamp 1676382929
transform 1 0 72000 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1332_
timestamp 1676382929
transform 1 0 72384 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1333_
timestamp 1676382929
transform 1 0 72768 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1334_
timestamp 1676382929
transform 1 0 73248 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1335_
timestamp 1676382929
transform 1 0 73632 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1336_
timestamp 1676382929
transform 1 0 74016 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1337_
timestamp 1676382929
transform 1 0 74400 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1338_
timestamp 1676382929
transform 1 0 74784 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1339_
timestamp 1676382929
transform 1 0 75168 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1340_
timestamp 1676382929
transform 1 0 75552 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1341_
timestamp 1676382929
transform 1 0 76032 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1342_
timestamp 1676382929
transform -1 0 77088 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1343_
timestamp 1676382929
transform -1 0 77376 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1344_
timestamp 1676382929
transform 1 0 77376 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1345_
timestamp 1676382929
transform 1 0 77664 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1346_
timestamp 1676382929
transform 1 0 78048 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1347_
timestamp 1676382929
transform 1 0 78432 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1348_
timestamp 1676382929
transform 1 0 78720 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1349_
timestamp 1676382929
transform 1 0 79104 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1350_
timestamp 1676382929
transform 1 0 78528 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1351_
timestamp 1676382929
transform 1 0 78144 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1352_
timestamp 1676382929
transform 1 0 77760 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1353_
timestamp 1676382929
transform 1 0 77376 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1354_
timestamp 1676382929
transform 1 0 77088 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1355_
timestamp 1676382929
transform -1 0 77088 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1356_
timestamp 1676382929
transform -1 0 76704 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1357_
timestamp 1676382929
transform 1 0 75648 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1358_
timestamp 1676382929
transform 1 0 75264 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1359_
timestamp 1676382929
transform 1 0 74880 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1360_
timestamp 1676382929
transform 1 0 74496 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1361_
timestamp 1676382929
transform 1 0 74112 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1362_
timestamp 1676382929
transform 1 0 73632 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1363_
timestamp 1676382929
transform 1 0 73248 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1364_
timestamp 1676382929
transform 1 0 72864 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1365_
timestamp 1676382929
transform 1 0 72480 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1366_
timestamp 1676382929
transform 1 0 72096 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1367_
timestamp 1676382929
transform 1 0 71712 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1368_
timestamp 1676382929
transform 1 0 71232 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1369_
timestamp 1676382929
transform 1 0 70848 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1370_
timestamp 1676382929
transform 1 0 70464 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1371_
timestamp 1676382929
transform 1 0 70080 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1372_
timestamp 1676382929
transform 1 0 69696 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1373_
timestamp 1676382929
transform 1 0 69312 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1374_
timestamp 1676382929
transform 1 0 68928 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1375_
timestamp 1676382929
transform 1 0 68448 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1376_
timestamp 1676382929
transform 1 0 68064 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1377_
timestamp 1676382929
transform 1 0 67680 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1378_
timestamp 1676382929
transform 1 0 67296 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1379_
timestamp 1676382929
transform 1 0 66912 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1380_
timestamp 1676382929
transform 1 0 66432 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1381_
timestamp 1676382929
transform 1 0 66048 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1382_
timestamp 1676382929
transform 1 0 65664 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1383_
timestamp 1676382929
transform 1 0 65280 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1384_
timestamp 1676382929
transform 1 0 64896 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1385_
timestamp 1676382929
transform 1 0 64416 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1386_
timestamp 1676382929
transform 1 0 64032 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1387_
timestamp 1676382929
transform 1 0 63744 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1388_
timestamp 1676382929
transform 1 0 63456 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1389_
timestamp 1676382929
transform 1 0 63168 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1390_
timestamp 1676382929
transform 1 0 62880 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1391_
timestamp 1676382929
transform 1 0 62592 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1392_
timestamp 1676382929
transform 1 0 62304 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1393_
timestamp 1676382929
transform 1 0 62016 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1394_
timestamp 1676382929
transform 1 0 61344 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1395_
timestamp 1676382929
transform 1 0 60480 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1396_
timestamp 1676382929
transform 1 0 60000 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1397_
timestamp 1676382929
transform 1 0 59616 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1398_
timestamp 1676382929
transform 1 0 59232 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1399_
timestamp 1676382929
transform 1 0 58848 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1400_
timestamp 1676382929
transform 1 0 58464 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1401_
timestamp 1676382929
transform 1 0 58176 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1402_
timestamp 1676382929
transform 1 0 57888 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1403_
timestamp 1676382929
transform 1 0 57216 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1404_
timestamp 1676382929
transform 1 0 56832 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1405_
timestamp 1676382929
transform 1 0 56448 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1406_
timestamp 1676382929
transform 1 0 56064 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1407_
timestamp 1676382929
transform 1 0 55584 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1408_
timestamp 1676382929
transform 1 0 55200 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1409_
timestamp 1676382929
transform 1 0 54720 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1410_
timestamp 1676382929
transform 1 0 54336 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1411_
timestamp 1676382929
transform 1 0 52224 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1412_
timestamp 1676382929
transform 1 0 52224 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1413_
timestamp 1676382929
transform 1 0 5376 0 1 20412
box -48 -56 336 834
use sg13g2_mux2_1  _1414_
timestamp 1677247768
transform 1 0 22560 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1415_
timestamp 1676557249
transform -1 0 23424 0 -1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1416_
timestamp 1676627187
transform -1 0 2208 0 -1 23436
box -48 -56 432 834
use sg13g2_or2_1  _1417_
timestamp 1684236171
transform 1 0 1344 0 -1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _1418_
timestamp 1683973020
transform -1 0 3456 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1419_
timestamp 1685175443
transform -1 0 23136 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1420_
timestamp 1683973020
transform -1 0 22752 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1421_
timestamp 1677247768
transform -1 0 27648 0 1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1422_
timestamp 1676557249
transform -1 0 26688 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1423_
timestamp 1683973020
transform -1 0 25728 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1424_
timestamp 1685175443
transform -1 0 26784 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1425_
timestamp 1683973020
transform -1 0 26304 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1426_
timestamp 1677247768
transform 1 0 30048 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1427_
timestamp 1676557249
transform 1 0 31008 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1428_
timestamp 1683973020
transform -1 0 29088 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1429_
timestamp 1685175443
transform -1 0 30048 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1430_
timestamp 1683973020
transform -1 0 29568 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1431_
timestamp 1677247768
transform -1 0 33792 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1432_
timestamp 1676557249
transform 1 0 33024 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1433_
timestamp 1683973020
transform -1 0 32256 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1434_
timestamp 1685175443
transform -1 0 33024 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1435_
timestamp 1683973020
transform -1 0 32544 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1436_
timestamp 1677247768
transform -1 0 36960 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1437_
timestamp 1676557249
transform -1 0 36000 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1438_
timestamp 1683973020
transform -1 0 35328 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1439_
timestamp 1685175443
transform -1 0 36384 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1440_
timestamp 1683973020
transform -1 0 35904 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1441_
timestamp 1677247768
transform -1 0 39936 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1442_
timestamp 1676557249
transform 1 0 37440 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1443_
timestamp 1683973020
transform -1 0 38304 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1444_
timestamp 1685175443
transform -1 0 39456 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1445_
timestamp 1683973020
transform -1 0 38688 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1446_
timestamp 1677247768
transform 1 0 42720 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1447_
timestamp 1676557249
transform 1 0 43488 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1448_
timestamp 1683973020
transform -1 0 41376 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1449_
timestamp 1685175443
transform -1 0 42624 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1450_
timestamp 1683973020
transform -1 0 42336 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1451_
timestamp 1677247768
transform 1 0 42048 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1452_
timestamp 1676557249
transform 1 0 43968 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1453_
timestamp 1683973020
transform 1 0 42336 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1454_
timestamp 1685175443
transform -1 0 42048 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1455_
timestamp 1683973020
transform 1 0 41856 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1456_
timestamp 1677247768
transform -1 0 43776 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1457_
timestamp 1676557249
transform -1 0 43008 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1458_
timestamp 1683973020
transform 1 0 41760 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1459_
timestamp 1685175443
transform 1 0 41184 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1460_
timestamp 1683973020
transform 1 0 41472 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1461_
timestamp 1677247768
transform -1 0 40320 0 -1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1462_
timestamp 1676557249
transform 1 0 38976 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1463_
timestamp 1683973020
transform -1 0 40224 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1464_
timestamp 1685175443
transform 1 0 39072 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1465_
timestamp 1683973020
transform 1 0 39936 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1466_
timestamp 1677247768
transform -1 0 37632 0 1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1467_
timestamp 1676557249
transform -1 0 36672 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1468_
timestamp 1683973020
transform 1 0 38208 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1469_
timestamp 1685175443
transform 1 0 35904 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1470_
timestamp 1683973020
transform 1 0 37440 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1471_
timestamp 1677247768
transform 1 0 33504 0 1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1472_
timestamp 1676557249
transform 1 0 34464 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1473_
timestamp 1683973020
transform 1 0 34368 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1474_
timestamp 1685175443
transform 1 0 33216 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1475_
timestamp 1683973020
transform 1 0 33696 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1476_
timestamp 1677247768
transform -1 0 32928 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1477_
timestamp 1676557249
transform 1 0 32256 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1478_
timestamp 1683973020
transform 1 0 32736 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1479_
timestamp 1685175443
transform -1 0 33120 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1480_
timestamp 1683973020
transform -1 0 33120 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1481_
timestamp 1677247768
transform -1 0 37344 0 -1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1482_
timestamp 1676557249
transform -1 0 36480 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1483_
timestamp 1683973020
transform -1 0 35232 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1484_
timestamp 1685175443
transform -1 0 35712 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1485_
timestamp 1683973020
transform 1 0 34752 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1486_
timestamp 1677247768
transform -1 0 39360 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1487_
timestamp 1676557249
transform -1 0 38400 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1488_
timestamp 1683973020
transform -1 0 36480 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1489_
timestamp 1685175443
transform -1 0 37248 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1490_
timestamp 1683973020
transform -1 0 36768 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1491_
timestamp 1677247768
transform 1 0 41376 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1492_
timestamp 1676557249
transform 1 0 42336 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1493_
timestamp 1683973020
transform -1 0 39552 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1494_
timestamp 1685175443
transform -1 0 40992 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1495_
timestamp 1683973020
transform -1 0 40320 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1496_
timestamp 1677247768
transform 1 0 43296 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1497_
timestamp 1676557249
transform 1 0 44256 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1498_
timestamp 1683973020
transform -1 0 42048 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1499_
timestamp 1685175443
transform -1 0 43008 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1500_
timestamp 1683973020
transform -1 0 42528 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1501_
timestamp 1677247768
transform -1 0 47136 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1502_
timestamp 1676557249
transform -1 0 46176 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1503_
timestamp 1683973020
transform -1 0 44544 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1504_
timestamp 1685175443
transform -1 0 45792 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1505_
timestamp 1683973020
transform -1 0 45216 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1506_
timestamp 1677247768
transform 1 0 47808 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1507_
timestamp 1676557249
transform -1 0 48768 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1508_
timestamp 1683973020
transform -1 0 47136 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1509_
timestamp 1685175443
transform -1 0 47616 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1510_
timestamp 1683973020
transform -1 0 47616 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1511_
timestamp 1677247768
transform 1 0 47904 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1512_
timestamp 1676557249
transform -1 0 48672 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1513_
timestamp 1683973020
transform 1 0 47616 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1514_
timestamp 1685175443
transform -1 0 47808 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1515_
timestamp 1683973020
transform 1 0 47136 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1516_
timestamp 1677247768
transform 1 0 51456 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1517_
timestamp 1676557249
transform 1 0 52416 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1518_
timestamp 1683973020
transform -1 0 49248 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1519_
timestamp 1685175443
transform -1 0 50976 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1520_
timestamp 1683973020
transform -1 0 50400 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1521_
timestamp 1677247768
transform 1 0 53664 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1522_
timestamp 1676557249
transform -1 0 54624 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1523_
timestamp 1683973020
transform -1 0 52416 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1524_
timestamp 1685175443
transform -1 0 53088 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1525_
timestamp 1683973020
transform -1 0 52608 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1526_
timestamp 1677247768
transform 1 0 53088 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1527_
timestamp 1676557249
transform -1 0 54048 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1528_
timestamp 1683973020
transform 1 0 53184 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1529_
timestamp 1685175443
transform -1 0 53472 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1530_
timestamp 1683973020
transform 1 0 52704 0 1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _1531_
timestamp 1677247768
transform 1 0 52512 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1532_
timestamp 1676557249
transform 1 0 53472 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1533_
timestamp 1683973020
transform 1 0 52608 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1534_
timestamp 1685175443
transform 1 0 52128 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1535_
timestamp 1683973020
transform 1 0 52896 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1536_
timestamp 1677247768
transform 1 0 50592 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1537_
timestamp 1676557249
transform -1 0 51648 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1538_
timestamp 1683973020
transform 1 0 51264 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1539_
timestamp 1685175443
transform 1 0 50112 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1540_
timestamp 1683973020
transform 1 0 50688 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1541_
timestamp 1677247768
transform 1 0 48000 0 -1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1542_
timestamp 1676557249
transform -1 0 48960 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1543_
timestamp 1683973020
transform 1 0 49056 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1544_
timestamp 1685175443
transform 1 0 47808 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1545_
timestamp 1683973020
transform 1 0 48192 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1546_
timestamp 1677247768
transform 1 0 46752 0 -1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1547_
timestamp 1676557249
transform -1 0 47712 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1548_
timestamp 1683973020
transform 1 0 47232 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1549_
timestamp 1685175443
transform 1 0 46272 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1550_
timestamp 1683973020
transform 1 0 46752 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1551_
timestamp 1677247768
transform 1 0 45216 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1552_
timestamp 1676557249
transform 1 0 46272 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1553_
timestamp 1683973020
transform 1 0 45504 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1554_
timestamp 1685175443
transform -1 0 45792 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1555_
timestamp 1683973020
transform 1 0 45792 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1556_
timestamp 1677247768
transform -1 0 49248 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1557_
timestamp 1676557249
transform -1 0 48288 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1558_
timestamp 1683973020
transform -1 0 46464 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1559_
timestamp 1685175443
transform -1 0 47808 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1560_
timestamp 1683973020
transform -1 0 47136 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1561_
timestamp 1677247768
transform 1 0 50208 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1562_
timestamp 1676557249
transform 1 0 51168 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1563_
timestamp 1683973020
transform -1 0 49056 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1564_
timestamp 1685175443
transform -1 0 50112 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1565_
timestamp 1683973020
transform -1 0 49536 0 -1 17388
box -48 -56 528 834
use sg13g2_mux2_1  _1566_
timestamp 1677247768
transform 1 0 52032 0 -1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1567_
timestamp 1676557249
transform 1 0 52800 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1568_
timestamp 1683973020
transform -1 0 51264 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1569_
timestamp 1685175443
transform -1 0 51936 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1570_
timestamp 1683973020
transform -1 0 51552 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1571_
timestamp 1677247768
transform 1 0 55872 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1572_
timestamp 1676557249
transform -1 0 56736 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1573_
timestamp 1683973020
transform -1 0 53760 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1574_
timestamp 1685175443
transform -1 0 55488 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1575_
timestamp 1683973020
transform -1 0 54816 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1576_
timestamp 1677247768
transform 1 0 57696 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1577_
timestamp 1676557249
transform -1 0 58560 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1578_
timestamp 1683973020
transform -1 0 56448 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1579_
timestamp 1685175443
transform -1 0 56928 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1580_
timestamp 1683973020
transform 1 0 56448 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1581_
timestamp 1677247768
transform -1 0 59904 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1582_
timestamp 1676557249
transform 1 0 59040 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1583_
timestamp 1683973020
transform 1 0 57600 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1584_
timestamp 1685175443
transform -1 0 58560 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1585_
timestamp 1683973020
transform -1 0 58176 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1586_
timestamp 1677247768
transform 1 0 58176 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1587_
timestamp 1676557249
transform 1 0 59520 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1588_
timestamp 1683973020
transform 1 0 58176 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1589_
timestamp 1685175443
transform -1 0 58176 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1590_
timestamp 1683973020
transform 1 0 57696 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1591_
timestamp 1677247768
transform 1 0 59520 0 1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1592_
timestamp 1676557249
transform -1 0 60480 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1593_
timestamp 1683973020
transform -1 0 58944 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1594_
timestamp 1685175443
transform -1 0 58944 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1595_
timestamp 1683973020
transform 1 0 57984 0 -1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _1596_
timestamp 1677247768
transform 1 0 60192 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1597_
timestamp 1676557249
transform 1 0 61344 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1598_
timestamp 1683973020
transform -1 0 59616 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1599_
timestamp 1685175443
transform 1 0 58848 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1600_
timestamp 1683973020
transform 1 0 59136 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1601_
timestamp 1677247768
transform 1 0 55968 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1602_
timestamp 1676557249
transform -1 0 56928 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1603_
timestamp 1683973020
transform 1 0 57888 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1604_
timestamp 1685175443
transform -1 0 55968 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1605_
timestamp 1683973020
transform 1 0 56928 0 1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1606_
timestamp 1677247768
transform 1 0 55968 0 1 756
box -48 -56 1008 834
use sg13g2_nand2_1  _1607_
timestamp 1676557249
transform -1 0 57120 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1608_
timestamp 1683973020
transform -1 0 56160 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1609_
timestamp 1685175443
transform -1 0 55872 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1610_
timestamp 1683973020
transform 1 0 55968 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1611_
timestamp 1677247768
transform 1 0 59232 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1612_
timestamp 1676557249
transform 1 0 60192 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1613_
timestamp 1683973020
transform -1 0 57600 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1614_
timestamp 1685175443
transform -1 0 60768 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1615_
timestamp 1683973020
transform -1 0 59040 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1616_
timestamp 1677247768
transform 1 0 63648 0 1 756
box -48 -56 1008 834
use sg13g2_nand2_1  _1617_
timestamp 1676557249
transform 1 0 64608 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _1618_
timestamp 1683973020
transform -1 0 62112 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _1619_
timestamp 1685175443
transform -1 0 63072 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1620_
timestamp 1683973020
transform -1 0 62592 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1621_
timestamp 1677247768
transform 1 0 65376 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1622_
timestamp 1676557249
transform -1 0 66432 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1623_
timestamp 1683973020
transform -1 0 64128 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1624_
timestamp 1685175443
transform -1 0 64704 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1625_
timestamp 1683973020
transform -1 0 64224 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1626_
timestamp 1677247768
transform 1 0 65472 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1627_
timestamp 1676557249
transform -1 0 66528 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1628_
timestamp 1683973020
transform 1 0 65472 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1629_
timestamp 1685175443
transform -1 0 65472 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1630_
timestamp 1683973020
transform 1 0 64512 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1631_
timestamp 1677247768
transform 1 0 64512 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1632_
timestamp 1676557249
transform -1 0 65568 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1633_
timestamp 1683973020
transform 1 0 64704 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1634_
timestamp 1685175443
transform -1 0 64512 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1635_
timestamp 1683973020
transform 1 0 63552 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1636_
timestamp 1677247768
transform 1 0 64128 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1637_
timestamp 1676557249
transform -1 0 64896 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1638_
timestamp 1683973020
transform 1 0 64224 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1639_
timestamp 1685175443
transform 1 0 63744 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1640_
timestamp 1683973020
transform 1 0 64704 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1641_
timestamp 1677247768
transform 1 0 63264 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1642_
timestamp 1676557249
transform -1 0 64224 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1643_
timestamp 1683973020
transform 1 0 63360 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1644_
timestamp 1685175443
transform 1 0 62688 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1645_
timestamp 1683973020
transform 1 0 62976 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1646_
timestamp 1677247768
transform -1 0 61920 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1647_
timestamp 1676557249
transform -1 0 61152 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1648_
timestamp 1683973020
transform 1 0 62016 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1649_
timestamp 1685175443
transform -1 0 62400 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1650_
timestamp 1683973020
transform 1 0 61248 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1651_
timestamp 1677247768
transform -1 0 64992 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1652_
timestamp 1676557249
transform -1 0 64032 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1653_
timestamp 1683973020
transform -1 0 64224 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1654_
timestamp 1685175443
transform -1 0 64224 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1655_
timestamp 1683973020
transform -1 0 64704 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1656_
timestamp 1677247768
transform 1 0 69504 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1657_
timestamp 1676557249
transform -1 0 70368 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1658_
timestamp 1683973020
transform -1 0 67680 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1659_
timestamp 1685175443
transform -1 0 68928 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1660_
timestamp 1683973020
transform -1 0 68448 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1661_
timestamp 1677247768
transform -1 0 70368 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1662_
timestamp 1676557249
transform -1 0 69984 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1663_
timestamp 1683973020
transform 1 0 69024 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1664_
timestamp 1685175443
transform -1 0 69024 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1665_
timestamp 1683973020
transform 1 0 68832 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1666_
timestamp 1677247768
transform 1 0 69120 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1667_
timestamp 1676557249
transform -1 0 69984 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1668_
timestamp 1683973020
transform 1 0 68928 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1669_
timestamp 1685175443
transform -1 0 68640 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1670_
timestamp 1683973020
transform 1 0 68640 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1671_
timestamp 1677247768
transform 1 0 70656 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1672_
timestamp 1676557249
transform -1 0 71616 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1673_
timestamp 1683973020
transform 1 0 69120 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1674_
timestamp 1685175443
transform -1 0 69984 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1675_
timestamp 1683973020
transform 1 0 68640 0 1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1676_
timestamp 1677247768
transform 1 0 71136 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1677_
timestamp 1676557249
transform 1 0 72096 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1678_
timestamp 1683973020
transform 1 0 69984 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1679_
timestamp 1685175443
transform 1 0 69216 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1680_
timestamp 1683973020
transform 1 0 69696 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1681_
timestamp 1677247768
transform 1 0 67776 0 -1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1682_
timestamp 1676557249
transform 1 0 68544 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1683_
timestamp 1683973020
transform 1 0 68736 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1684_
timestamp 1685175443
transform -1 0 68544 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1685_
timestamp 1683973020
transform 1 0 67296 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1686_
timestamp 1677247768
transform -1 0 72000 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1687_
timestamp 1676557249
transform 1 0 71136 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1688_
timestamp 1683973020
transform -1 0 69024 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1689_
timestamp 1685175443
transform -1 0 70080 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1690_
timestamp 1683973020
transform -1 0 69504 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1691_
timestamp 1677247768
transform -1 0 74208 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1692_
timestamp 1676557249
transform -1 0 73152 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1693_
timestamp 1683973020
transform -1 0 71040 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1694_
timestamp 1685175443
transform -1 0 72000 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1695_
timestamp 1683973020
transform -1 0 71520 0 1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1696_
timestamp 1677247768
transform 1 0 76608 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1697_
timestamp 1676557249
transform 1 0 77568 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1698_
timestamp 1683973020
transform -1 0 74976 0 -1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1699_
timestamp 1685175443
transform -1 0 76320 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1700_
timestamp 1683973020
transform -1 0 75552 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1701_
timestamp 1677247768
transform 1 0 76224 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1702_
timestamp 1676557249
transform 1 0 77184 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1703_
timestamp 1683973020
transform 1 0 76128 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1704_
timestamp 1685175443
transform 1 0 75744 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1705_
timestamp 1683973020
transform 1 0 76320 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1706_
timestamp 1677247768
transform 1 0 76032 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1707_
timestamp 1676557249
transform 1 0 76896 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1708_
timestamp 1683973020
transform -1 0 76320 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1709_
timestamp 1685175443
transform 1 0 75552 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1710_
timestamp 1683973020
transform 1 0 76128 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1711_
timestamp 1677247768
transform 1 0 76032 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1712_
timestamp 1676557249
transform -1 0 76896 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1713_
timestamp 1683973020
transform 1 0 75936 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1714_
timestamp 1685175443
transform -1 0 76512 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1715_
timestamp 1683973020
transform 1 0 75456 0 1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _1716_
timestamp 1677247768
transform 1 0 76032 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1717_
timestamp 1676557249
transform 1 0 76992 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1718_
timestamp 1683973020
transform 1 0 75552 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1719_
timestamp 1685175443
transform -1 0 75936 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1720_
timestamp 1683973020
transform 1 0 75936 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1721_
timestamp 1677247768
transform 1 0 75168 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1722_
timestamp 1676557249
transform 1 0 76032 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1723_
timestamp 1683973020
transform 1 0 75552 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1724_
timestamp 1685175443
transform -1 0 75072 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1725_
timestamp 1683973020
transform 1 0 75072 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1726_
timestamp 1677247768
transform 1 0 75264 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1727_
timestamp 1676557249
transform -1 0 76320 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1728_
timestamp 1683973020
transform 1 0 74688 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1729_
timestamp 1685175443
transform -1 0 75168 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1730_
timestamp 1683973020
transform 1 0 74208 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1731_
timestamp 1677247768
transform 1 0 74496 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1732_
timestamp 1676557249
transform -1 0 75456 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1733_
timestamp 1683973020
transform 1 0 74688 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1734_
timestamp 1685175443
transform -1 0 74496 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1735_
timestamp 1683973020
transform 1 0 73536 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1736_
timestamp 1677247768
transform 1 0 75264 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1737_
timestamp 1676557249
transform -1 0 76128 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1738_
timestamp 1683973020
transform 1 0 74208 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1739_
timestamp 1685175443
transform -1 0 75072 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1740_
timestamp 1683973020
transform -1 0 74592 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1741_
timestamp 1677247768
transform 1 0 76032 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1742_
timestamp 1676557249
transform -1 0 76992 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1743_
timestamp 1683973020
transform 1 0 75072 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1744_
timestamp 1685175443
transform -1 0 76032 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1745_
timestamp 1683973020
transform 1 0 74784 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1746_
timestamp 1677247768
transform 1 0 75936 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1747_
timestamp 1676557249
transform -1 0 76800 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1748_
timestamp 1683973020
transform 1 0 75360 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1749_
timestamp 1685175443
transform -1 0 75648 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1750_
timestamp 1683973020
transform 1 0 75168 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1751_
timestamp 1677247768
transform 1 0 76032 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1752_
timestamp 1676557249
transform 1 0 76896 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1753_
timestamp 1683973020
transform 1 0 75648 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1754_
timestamp 1685175443
transform -1 0 75264 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1755_
timestamp 1683973020
transform 1 0 75264 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1756_
timestamp 1677247768
transform 1 0 77280 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1757_
timestamp 1676557249
transform -1 0 78624 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1758_
timestamp 1683973020
transform 1 0 75744 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1759_
timestamp 1685175443
transform -1 0 76608 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1760_
timestamp 1683973020
transform -1 0 76128 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1761_
timestamp 1677247768
transform 1 0 76416 0 1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1762_
timestamp 1676557249
transform -1 0 77376 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1763_
timestamp 1683973020
transform 1 0 76608 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1764_
timestamp 1685175443
transform -1 0 76416 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1765_
timestamp 1683973020
transform 1 0 75936 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1766_
timestamp 1677247768
transform 1 0 76704 0 -1 38556
box -48 -56 1008 834
use sg13g2_nand2_1  _1767_
timestamp 1676557249
transform -1 0 77760 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1768_
timestamp 1683973020
transform 1 0 76416 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1769_
timestamp 1685175443
transform 1 0 74976 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1770_
timestamp 1683973020
transform 1 0 76032 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1771_
timestamp 1677247768
transform 1 0 72576 0 1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1772_
timestamp 1676557249
transform 1 0 73920 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1773_
timestamp 1683973020
transform 1 0 74208 0 1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1774_
timestamp 1685175443
transform 1 0 72672 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1775_
timestamp 1683973020
transform 1 0 73632 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1776_
timestamp 1677247768
transform 1 0 70848 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1777_
timestamp 1676557249
transform 1 0 72288 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1778_
timestamp 1683973020
transform 1 0 71808 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1779_
timestamp 1685175443
transform 1 0 70368 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1780_
timestamp 1683973020
transform 1 0 71808 0 -1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _1781_
timestamp 1677247768
transform 1 0 67872 0 1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1782_
timestamp 1676557249
transform 1 0 68832 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _1783_
timestamp 1683973020
transform 1 0 69600 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1784_
timestamp 1685175443
transform 1 0 67968 0 -1 38556
box -48 -56 538 834
use sg13g2_a21oi_1  _1785_
timestamp 1683973020
transform 1 0 68352 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1786_
timestamp 1677247768
transform 1 0 66240 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1787_
timestamp 1676557249
transform -1 0 67584 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1788_
timestamp 1683973020
transform 1 0 67008 0 1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1789_
timestamp 1685175443
transform -1 0 66240 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1790_
timestamp 1683973020
transform 1 0 66720 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _1791_
timestamp 1677247768
transform -1 0 66624 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1792_
timestamp 1676557249
transform -1 0 65664 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1793_
timestamp 1683973020
transform 1 0 66048 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1794_
timestamp 1685175443
transform 1 0 65952 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1795_
timestamp 1683973020
transform 1 0 66432 0 1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _1796_
timestamp 1677247768
transform 1 0 71424 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1797_
timestamp 1676557249
transform 1 0 72384 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1798_
timestamp 1683973020
transform -1 0 69216 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1799_
timestamp 1685175443
transform -1 0 70656 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1800_
timestamp 1683973020
transform -1 0 70176 0 -1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _1801_
timestamp 1677247768
transform 1 0 70752 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1802_
timestamp 1676557249
transform -1 0 71712 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1803_
timestamp 1683973020
transform -1 0 71232 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1804_
timestamp 1685175443
transform -1 0 70848 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1805_
timestamp 1683973020
transform 1 0 70752 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1806_
timestamp 1677247768
transform 1 0 70080 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1807_
timestamp 1676557249
transform -1 0 70944 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1808_
timestamp 1683973020
transform 1 0 70272 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1809_
timestamp 1685175443
transform -1 0 70656 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1810_
timestamp 1683973020
transform 1 0 69792 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1811_
timestamp 1677247768
transform 1 0 70752 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1812_
timestamp 1676557249
transform 1 0 71712 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1813_
timestamp 1683973020
transform 1 0 69984 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1814_
timestamp 1685175443
transform 1 0 69216 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1815_
timestamp 1683973020
transform 1 0 69504 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1816_
timestamp 1677247768
transform 1 0 66912 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1817_
timestamp 1676557249
transform -1 0 68448 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1818_
timestamp 1683973020
transform 1 0 68256 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1819_
timestamp 1685175443
transform 1 0 67104 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1820_
timestamp 1683973020
transform 1 0 67584 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1821_
timestamp 1677247768
transform 1 0 62976 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1822_
timestamp 1676557249
transform -1 0 63840 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1823_
timestamp 1683973020
transform 1 0 65280 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1824_
timestamp 1685175443
transform 1 0 64128 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1825_
timestamp 1683973020
transform 1 0 64608 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1826_
timestamp 1677247768
transform -1 0 65376 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1827_
timestamp 1676557249
transform 1 0 64704 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1828_
timestamp 1683973020
transform 1 0 63744 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1829_
timestamp 1685175443
transform 1 0 63744 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1830_
timestamp 1683973020
transform -1 0 64128 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1831_
timestamp 1677247768
transform -1 0 65952 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1832_
timestamp 1676557249
transform -1 0 64992 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1833_
timestamp 1683973020
transform 1 0 63264 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1834_
timestamp 1685175443
transform 1 0 63168 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1835_
timestamp 1683973020
transform 1 0 63648 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1836_
timestamp 1677247768
transform 1 0 62880 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1837_
timestamp 1676557249
transform 1 0 63840 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1838_
timestamp 1683973020
transform 1 0 62592 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1839_
timestamp 1685175443
transform -1 0 62784 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1840_
timestamp 1683973020
transform 1 0 62496 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1841_
timestamp 1677247768
transform -1 0 63264 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1842_
timestamp 1676557249
transform 1 0 62592 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1843_
timestamp 1683973020
transform 1 0 62112 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1844_
timestamp 1685175443
transform -1 0 62208 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1845_
timestamp 1683973020
transform 1 0 61824 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1846_
timestamp 1677247768
transform 1 0 62976 0 -1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1847_
timestamp 1676557249
transform 1 0 63936 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _1848_
timestamp 1683973020
transform 1 0 61248 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1849_
timestamp 1685175443
transform 1 0 61344 0 -1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1850_
timestamp 1683973020
transform 1 0 61824 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1851_
timestamp 1677247768
transform 1 0 58080 0 -1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1852_
timestamp 1676557249
transform 1 0 58752 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1853_
timestamp 1683973020
transform 1 0 60096 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1854_
timestamp 1685175443
transform 1 0 58464 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1855_
timestamp 1683973020
transform 1 0 57984 0 -1 38556
box -48 -56 528 834
use sg13g2_mux2_1  _1856_
timestamp 1677247768
transform -1 0 56448 0 1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1857_
timestamp 1676557249
transform -1 0 55008 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1858_
timestamp 1683973020
transform 1 0 56928 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1859_
timestamp 1685175443
transform -1 0 56160 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1860_
timestamp 1683973020
transform 1 0 55392 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1861_
timestamp 1677247768
transform 1 0 58176 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1862_
timestamp 1676557249
transform 1 0 59136 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1863_
timestamp 1683973020
transform 1 0 58080 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1864_
timestamp 1685175443
transform -1 0 58752 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1865_
timestamp 1683973020
transform -1 0 57888 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1866_
timestamp 1677247768
transform 1 0 59616 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1867_
timestamp 1676557249
transform 1 0 60768 0 -1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1868_
timestamp 1683973020
transform -1 0 60000 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1869_
timestamp 1685175443
transform -1 0 59616 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1870_
timestamp 1683973020
transform 1 0 59520 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1871_
timestamp 1677247768
transform 1 0 59328 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1872_
timestamp 1676557249
transform 1 0 60576 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1873_
timestamp 1683973020
transform -1 0 60000 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1874_
timestamp 1685175443
transform 1 0 59040 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1875_
timestamp 1683973020
transform 1 0 59808 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1876_
timestamp 1677247768
transform -1 0 60000 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1877_
timestamp 1676557249
transform -1 0 59616 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1878_
timestamp 1683973020
transform 1 0 58752 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1879_
timestamp 1685175443
transform 1 0 57984 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1880_
timestamp 1683973020
transform 1 0 58272 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1881_
timestamp 1677247768
transform -1 0 56256 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1882_
timestamp 1676557249
transform -1 0 55296 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1883_
timestamp 1683973020
transform 1 0 56736 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1884_
timestamp 1685175443
transform 1 0 55584 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1885_
timestamp 1683973020
transform 1 0 56256 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1886_
timestamp 1677247768
transform 1 0 55200 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1887_
timestamp 1676557249
transform -1 0 55968 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1888_
timestamp 1683973020
transform 1 0 55104 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1889_
timestamp 1685175443
transform -1 0 55872 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1890_
timestamp 1683973020
transform 1 0 54528 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1891_
timestamp 1677247768
transform 1 0 54912 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1892_
timestamp 1676557249
transform -1 0 55872 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1893_
timestamp 1683973020
transform 1 0 54720 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1894_
timestamp 1685175443
transform -1 0 55008 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1895_
timestamp 1683973020
transform 1 0 54432 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1896_
timestamp 1677247768
transform 1 0 54720 0 -1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1897_
timestamp 1676557249
transform -1 0 55296 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1898_
timestamp 1683973020
transform 1 0 54048 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1899_
timestamp 1685175443
transform 1 0 53568 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1900_
timestamp 1683973020
transform 1 0 53856 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1901_
timestamp 1677247768
transform -1 0 51936 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1902_
timestamp 1676557249
transform 1 0 51168 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1903_
timestamp 1683973020
transform 1 0 52128 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1904_
timestamp 1685175443
transform 1 0 50400 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1905_
timestamp 1683973020
transform 1 0 50880 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1906_
timestamp 1677247768
transform 1 0 46080 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1907_
timestamp 1676557249
transform -1 0 47808 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1908_
timestamp 1683973020
transform 1 0 49152 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1909_
timestamp 1685175443
transform -1 0 46848 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1910_
timestamp 1683973020
transform 1 0 46464 0 -1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _1911_
timestamp 1677247768
transform 1 0 50112 0 1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1912_
timestamp 1676557249
transform -1 0 51168 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1913_
timestamp 1683973020
transform -1 0 48960 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1914_
timestamp 1685175443
transform -1 0 49152 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1915_
timestamp 1683973020
transform 1 0 48864 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1916_
timestamp 1677247768
transform 1 0 50112 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1917_
timestamp 1676557249
transform -1 0 51072 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1918_
timestamp 1683973020
transform 1 0 49632 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1919_
timestamp 1685175443
transform -1 0 50112 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1920_
timestamp 1683973020
transform 1 0 49152 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1921_
timestamp 1677247768
transform 1 0 50976 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1922_
timestamp 1676557249
transform -1 0 51936 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1923_
timestamp 1683973020
transform 1 0 50112 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1924_
timestamp 1685175443
transform -1 0 50880 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1925_
timestamp 1683973020
transform 1 0 49920 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1926_
timestamp 1677247768
transform -1 0 52320 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1927_
timestamp 1676557249
transform -1 0 51360 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1928_
timestamp 1683973020
transform 1 0 50496 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1929_
timestamp 1685175443
transform 1 0 50496 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1930_
timestamp 1683973020
transform 1 0 51360 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1931_
timestamp 1677247768
transform 1 0 50112 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1932_
timestamp 1676557249
transform 1 0 51072 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1933_
timestamp 1683973020
transform 1 0 50304 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1934_
timestamp 1685175443
transform 1 0 49632 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1935_
timestamp 1683973020
transform 1 0 50496 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1936_
timestamp 1677247768
transform -1 0 50784 0 -1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _1937_
timestamp 1676557249
transform -1 0 49824 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _1938_
timestamp 1683973020
transform 1 0 49344 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1939_
timestamp 1685175443
transform 1 0 48480 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1940_
timestamp 1683973020
transform 1 0 48768 0 -1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1941_
timestamp 1677247768
transform 1 0 44832 0 -1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _1942_
timestamp 1676557249
transform 1 0 45888 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1943_
timestamp 1683973020
transform 1 0 46272 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1944_
timestamp 1685175443
transform 1 0 44736 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1945_
timestamp 1683973020
transform 1 0 45024 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1946_
timestamp 1677247768
transform 1 0 44928 0 1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1947_
timestamp 1676557249
transform 1 0 45888 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1948_
timestamp 1683973020
transform 1 0 44544 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1949_
timestamp 1685175443
transform -1 0 44352 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1950_
timestamp 1683973020
transform 1 0 44352 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1951_
timestamp 1677247768
transform -1 0 47040 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1952_
timestamp 1676557249
transform 1 0 46176 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1953_
timestamp 1683973020
transform 1 0 44832 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1954_
timestamp 1685175443
transform -1 0 44928 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1955_
timestamp 1683973020
transform 1 0 43968 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _1956_
timestamp 1677247768
transform 1 0 46080 0 -1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1957_
timestamp 1676557249
transform -1 0 46944 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1958_
timestamp 1683973020
transform 1 0 46368 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1959_
timestamp 1685175443
transform 1 0 45024 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1960_
timestamp 1683973020
transform 1 0 45504 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1961_
timestamp 1677247768
transform -1 0 46560 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1962_
timestamp 1676557249
transform 1 0 45792 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1963_
timestamp 1683973020
transform 1 0 44544 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1964_
timestamp 1685175443
transform 1 0 44832 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1965_
timestamp 1683973020
transform 1 0 45024 0 -1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1966_
timestamp 1677247768
transform -1 0 43584 0 1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1967_
timestamp 1676557249
transform 1 0 42816 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1968_
timestamp 1683973020
transform 1 0 43872 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1969_
timestamp 1685175443
transform 1 0 42336 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1970_
timestamp 1683973020
transform 1 0 42720 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1971_
timestamp 1677247768
transform -1 0 41952 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1972_
timestamp 1676557249
transform 1 0 41184 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1973_
timestamp 1683973020
transform 1 0 41568 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1974_
timestamp 1685175443
transform 1 0 40704 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1975_
timestamp 1683973020
transform 1 0 40992 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1976_
timestamp 1677247768
transform 1 0 40320 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1977_
timestamp 1676557249
transform -1 0 41376 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1978_
timestamp 1683973020
transform 1 0 40224 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1979_
timestamp 1685175443
transform 1 0 39840 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1980_
timestamp 1683973020
transform 1 0 40320 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1981_
timestamp 1677247768
transform 1 0 39360 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1982_
timestamp 1676557249
transform 1 0 40224 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1983_
timestamp 1683973020
transform 1 0 39648 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1984_
timestamp 1685175443
transform 1 0 39744 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1985_
timestamp 1683973020
transform 1 0 39168 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1986_
timestamp 1677247768
transform -1 0 41952 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1987_
timestamp 1676557249
transform -1 0 40800 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1988_
timestamp 1683973020
transform 1 0 39264 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1989_
timestamp 1685175443
transform 1 0 38784 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1990_
timestamp 1683973020
transform 1 0 38976 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1991_
timestamp 1677247768
transform 1 0 36096 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1992_
timestamp 1676557249
transform 1 0 37056 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1993_
timestamp 1683973020
transform 1 0 37728 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1994_
timestamp 1685175443
transform -1 0 36096 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1995_
timestamp 1683973020
transform 1 0 35808 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1996_
timestamp 1677247768
transform 1 0 34464 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1997_
timestamp 1676557249
transform -1 0 35328 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1998_
timestamp 1683973020
transform 1 0 35616 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1999_
timestamp 1685175443
transform 1 0 34176 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _2000_
timestamp 1683973020
transform 1 0 34656 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _2001_
timestamp 1677247768
transform 1 0 31872 0 1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _2002_
timestamp 1676557249
transform -1 0 32640 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2003_
timestamp 1683973020
transform 1 0 33120 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _2004_
timestamp 1685175443
transform 1 0 31872 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _2005_
timestamp 1683973020
transform 1 0 32352 0 -1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _2006_
timestamp 1677247768
transform 1 0 30720 0 1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _2007_
timestamp 1676557249
transform -1 0 31776 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2008_
timestamp 1683973020
transform 1 0 31104 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _2009_
timestamp 1685175443
transform 1 0 30240 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _2010_
timestamp 1683973020
transform 1 0 30624 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _2011_
timestamp 1677247768
transform 1 0 27744 0 -1 20412
box -48 -56 1008 834
use sg13g2_nand2_1  _2012_
timestamp 1676557249
transform 1 0 28704 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _2013_
timestamp 1683973020
transform 1 0 29280 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _2014_
timestamp 1685175443
transform 1 0 27744 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _2015_
timestamp 1683973020
transform 1 0 28224 0 -1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _2016_
timestamp 1677247768
transform 1 0 7488 0 1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _2017_
timestamp 1676557249
transform 1 0 8448 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2018_
timestamp 1683973020
transform 1 0 26592 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _2019_
timestamp 1685175443
transform 1 0 8448 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _2020_
timestamp 1683973020
transform 1 0 8256 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _2021_
timestamp 1677247768
transform 1 0 3360 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _2022_
timestamp 1676557249
transform 1 0 4224 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2023_
timestamp 1683973020
transform 1 0 2976 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _2024_
timestamp 1685175443
transform 1 0 2400 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _2025_
timestamp 1683973020
transform 1 0 2784 0 1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _2026_
timestamp 1677247768
transform -1 0 4704 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _2027_
timestamp 1676557249
transform -1 0 3744 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2028_
timestamp 1683973020
transform 1 0 2304 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _2029_
timestamp 1685175443
transform 1 0 1536 0 -1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _2030_
timestamp 1683973020
transform 1 0 2016 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _2031_
timestamp 1677247768
transform 1 0 3264 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _2032_
timestamp 1676557249
transform 1 0 4128 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2033_
timestamp 1683973020
transform 1 0 2496 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _2034_
timestamp 1685175443
transform 1 0 1728 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _2035_
timestamp 1683973020
transform 1 0 2016 0 -1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _2036_
timestamp 1677247768
transform 1 0 2688 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _2037_
timestamp 1676557249
transform 1 0 3648 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2038_
timestamp 1683973020
transform 1 0 2688 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _2039_
timestamp 1685175443
transform 1 0 1920 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _2040_
timestamp 1683973020
transform 1 0 2208 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _2041_
timestamp 1677247768
transform 1 0 3168 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _2042_
timestamp 1676557249
transform 1 0 4032 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2043_
timestamp 1683973020
transform 1 0 2592 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _2044_
timestamp 1685175443
transform 1 0 1920 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _2045_
timestamp 1683973020
transform 1 0 2112 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _2046_
timestamp 1677247768
transform 1 0 3840 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _2047_
timestamp 1676557249
transform 1 0 6528 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2048_
timestamp 1683973020
transform 1 0 2304 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _2049_
timestamp 1685175443
transform -1 0 2304 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _2050_
timestamp 1683973020
transform -1 0 2016 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _2051_
timestamp 1677247768
transform 1 0 2400 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _2052_
timestamp 1676557249
transform 1 0 3264 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2053_
timestamp 1683973020
transform 1 0 2688 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _2054_
timestamp 1685175443
transform 1 0 1440 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _2055_
timestamp 1683973020
transform 1 0 1920 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2056_
timestamp 1676557249
transform 1 0 22656 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2057_
timestamp 1683973020
transform 1 0 22560 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2058_
timestamp 1676557249
transform -1 0 27648 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2059_
timestamp 1683973020
transform 1 0 26688 0 -1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2060_
timestamp 1676557249
transform 1 0 30432 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2061_
timestamp 1683973020
transform 1 0 29856 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2062_
timestamp 1676557249
transform -1 0 33600 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2063_
timestamp 1683973020
transform 1 0 32448 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2064_
timestamp 1676557249
transform -1 0 36672 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2065_
timestamp 1683973020
transform 1 0 35616 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2066_
timestamp 1676557249
transform -1 0 38496 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2067_
timestamp 1683973020
transform -1 0 38976 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2068_
timestamp 1676557249
transform -1 0 44736 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2069_
timestamp 1683973020
transform 1 0 43872 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2070_
timestamp 1676557249
transform 1 0 42816 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2071_
timestamp 1683973020
transform 1 0 42624 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2072_
timestamp 1676557249
transform -1 0 43584 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2073_
timestamp 1683973020
transform 1 0 42720 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2074_
timestamp 1676557249
transform 1 0 39840 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2075_
timestamp 1683973020
transform 1 0 40320 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2076_
timestamp 1676557249
transform -1 0 37248 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2077_
timestamp 1683973020
transform -1 0 38112 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2078_
timestamp 1676557249
transform -1 0 34464 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2079_
timestamp 1683973020
transform 1 0 33696 0 -1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2080_
timestamp 1676557249
transform -1 0 32256 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2081_
timestamp 1683973020
transform 1 0 31392 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2082_
timestamp 1676557249
transform -1 0 36864 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2083_
timestamp 1683973020
transform -1 0 36960 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2084_
timestamp 1676557249
transform -1 0 39264 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2085_
timestamp 1683973020
transform 1 0 39360 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2086_
timestamp 1676557249
transform -1 0 42528 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2087_
timestamp 1683973020
transform -1 0 42240 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2088_
timestamp 1676557249
transform -1 0 43584 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2089_
timestamp 1683973020
transform -1 0 44064 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2090_
timestamp 1676557249
transform -1 0 47232 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2091_
timestamp 1683973020
transform 1 0 46176 0 1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2092_
timestamp 1676557249
transform -1 0 50016 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2093_
timestamp 1683973020
transform 1 0 48768 0 1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2094_
timestamp 1676557249
transform 1 0 48384 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2095_
timestamp 1683973020
transform 1 0 48864 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2096_
timestamp 1676557249
transform -1 0 52800 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2097_
timestamp 1683973020
transform 1 0 51456 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2098_
timestamp 1676557249
transform 1 0 54624 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2099_
timestamp 1683973020
transform 1 0 54048 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2100_
timestamp 1676557249
transform 1 0 54144 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2101_
timestamp 1683973020
transform 1 0 53952 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2102_
timestamp 1676557249
transform -1 0 54048 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2103_
timestamp 1683973020
transform 1 0 53280 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2104_
timestamp 1676557249
transform -1 0 51936 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2105_
timestamp 1683973020
transform -1 0 52032 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2106_
timestamp 1676557249
transform -1 0 49824 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2107_
timestamp 1683973020
transform 1 0 48960 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2108_
timestamp 1676557249
transform 1 0 47712 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2109_
timestamp 1683973020
transform 1 0 47520 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2110_
timestamp 1676557249
transform 1 0 46080 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2111_
timestamp 1683973020
transform 1 0 45888 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2112_
timestamp 1676557249
transform -1 0 49632 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2113_
timestamp 1683973020
transform 1 0 48960 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2114_
timestamp 1676557249
transform -1 0 51552 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2115_
timestamp 1683973020
transform -1 0 50208 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2116_
timestamp 1676557249
transform -1 0 53376 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2117_
timestamp 1683973020
transform 1 0 52512 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2118_
timestamp 1676557249
transform -1 0 57696 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2119_
timestamp 1683973020
transform 1 0 56832 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2120_
timestamp 1676557249
transform -1 0 58080 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2121_
timestamp 1683973020
transform 1 0 58656 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2122_
timestamp 1676557249
transform 1 0 59232 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2123_
timestamp 1683973020
transform 1 0 58752 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2124_
timestamp 1676557249
transform -1 0 60288 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2125_
timestamp 1683973020
transform 1 0 59040 0 1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2126_
timestamp 1676557249
transform 1 0 60000 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2127_
timestamp 1683973020
transform -1 0 60960 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2128_
timestamp 1676557249
transform -1 0 62112 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2129_
timestamp 1683973020
transform 1 0 60960 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2130_
timestamp 1676557249
transform -1 0 56544 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2131_
timestamp 1683973020
transform 1 0 55584 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2132_
timestamp 1676557249
transform -1 0 57312 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _2133_
timestamp 1683973020
transform 1 0 56256 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2134_
timestamp 1676557249
transform -1 0 59616 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2135_
timestamp 1683973020
transform 1 0 58752 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2136_
timestamp 1676557249
transform -1 0 64992 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2137_
timestamp 1683973020
transform 1 0 64128 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2138_
timestamp 1676557249
transform -1 0 66816 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2139_
timestamp 1683973020
transform 1 0 66048 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2140_
timestamp 1676557249
transform -1 0 66912 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2141_
timestamp 1683973020
transform 1 0 66240 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2142_
timestamp 1676557249
transform -1 0 66144 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2143_
timestamp 1683973020
transform 1 0 65472 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2144_
timestamp 1676557249
transform -1 0 65568 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2145_
timestamp 1683973020
transform 1 0 64896 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2146_
timestamp 1676557249
transform -1 0 64704 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2147_
timestamp 1683973020
transform -1 0 64704 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2148_
timestamp 1676557249
transform -1 0 62496 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2149_
timestamp 1683973020
transform 1 0 60864 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2150_
timestamp 1676557249
transform 1 0 64704 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2151_
timestamp 1683973020
transform -1 0 65472 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2152_
timestamp 1676557249
transform -1 0 71232 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2153_
timestamp 1683973020
transform -1 0 70464 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2154_
timestamp 1676557249
transform -1 0 70752 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2155_
timestamp 1683973020
transform -1 0 70368 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2156_
timestamp 1676557249
transform -1 0 71040 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2157_
timestamp 1683973020
transform 1 0 69792 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2158_
timestamp 1676557249
transform -1 0 72000 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2159_
timestamp 1683973020
transform 1 0 71328 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2160_
timestamp 1676557249
transform -1 0 72864 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2161_
timestamp 1683973020
transform 1 0 71616 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2162_
timestamp 1676557249
transform -1 0 69312 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2163_
timestamp 1683973020
transform -1 0 69024 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _2164_
timestamp 1676557249
transform -1 0 72384 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2165_
timestamp 1683973020
transform 1 0 71520 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2166_
timestamp 1676557249
transform 1 0 74208 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2167_
timestamp 1683973020
transform 1 0 73920 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2168_
timestamp 1676557249
transform -1 0 79008 0 -1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2169_
timestamp 1683973020
transform 1 0 78144 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2170_
timestamp 1676557249
transform -1 0 77952 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2171_
timestamp 1683973020
transform 1 0 77088 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2172_
timestamp 1676557249
transform -1 0 77760 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2173_
timestamp 1683973020
transform 1 0 77088 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2174_
timestamp 1676557249
transform -1 0 78240 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2175_
timestamp 1683973020
transform 1 0 76896 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2176_
timestamp 1676557249
transform -1 0 77856 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2177_
timestamp 1683973020
transform 1 0 76992 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2178_
timestamp 1676557249
transform -1 0 77184 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2179_
timestamp 1683973020
transform 1 0 76320 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2180_
timestamp 1676557249
transform -1 0 77280 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2181_
timestamp 1683973020
transform 1 0 76416 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2182_
timestamp 1676557249
transform -1 0 76128 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2183_
timestamp 1683973020
transform 1 0 75552 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2184_
timestamp 1676557249
transform -1 0 76800 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2185_
timestamp 1683973020
transform 1 0 76128 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2186_
timestamp 1676557249
transform -1 0 77472 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2187_
timestamp 1683973020
transform 1 0 76704 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2188_
timestamp 1676557249
transform -1 0 77568 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2189_
timestamp 1683973020
transform 1 0 76704 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2190_
timestamp 1676557249
transform -1 0 77760 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2191_
timestamp 1683973020
transform 1 0 76992 0 1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2192_
timestamp 1676557249
transform -1 0 76992 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2193_
timestamp 1683973020
transform 1 0 77184 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2194_
timestamp 1676557249
transform -1 0 78240 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2195_
timestamp 1683973020
transform 1 0 77376 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2196_
timestamp 1676557249
transform -1 0 78432 0 1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2197_
timestamp 1683973020
transform 1 0 76512 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2198_
timestamp 1676557249
transform -1 0 73920 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2199_
timestamp 1683973020
transform 1 0 73152 0 1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2200_
timestamp 1676557249
transform -1 0 71904 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2201_
timestamp 1683973020
transform -1 0 72096 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2202_
timestamp 1676557249
transform -1 0 69600 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2203_
timestamp 1683973020
transform -1 0 69120 0 -1 38556
box -48 -56 528 834
use sg13g2_nand2_1  _2204_
timestamp 1676557249
transform -1 0 67776 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2205_
timestamp 1683973020
transform 1 0 66912 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2206_
timestamp 1676557249
transform -1 0 67200 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2207_
timestamp 1683973020
transform 1 0 66336 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2208_
timestamp 1676557249
transform -1 0 72768 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2209_
timestamp 1683973020
transform 1 0 71904 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2210_
timestamp 1676557249
transform -1 0 72288 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _2211_
timestamp 1683973020
transform 1 0 71424 0 1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2212_
timestamp 1676557249
transform -1 0 71808 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2213_
timestamp 1683973020
transform 1 0 70944 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2214_
timestamp 1676557249
transform -1 0 71904 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2215_
timestamp 1683973020
transform 1 0 70656 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2216_
timestamp 1676557249
transform -1 0 68448 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2217_
timestamp 1683973020
transform 1 0 67584 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2218_
timestamp 1676557249
transform -1 0 64704 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2219_
timestamp 1683973020
transform 1 0 63840 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2220_
timestamp 1676557249
transform -1 0 65952 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2221_
timestamp 1683973020
transform 1 0 65088 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2222_
timestamp 1676557249
transform -1 0 66240 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2223_
timestamp 1683973020
transform 1 0 65568 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2224_
timestamp 1676557249
transform -1 0 64608 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2225_
timestamp 1683973020
transform 1 0 62976 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2226_
timestamp 1676557249
transform -1 0 63360 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2227_
timestamp 1683973020
transform 1 0 62496 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2228_
timestamp 1676557249
transform -1 0 64320 0 -1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _2229_
timestamp 1683973020
transform 1 0 63456 0 -1 38556
box -48 -56 528 834
use sg13g2_nand2_1  _2230_
timestamp 1676557249
transform -1 0 59904 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2231_
timestamp 1683973020
transform 1 0 59040 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2232_
timestamp 1676557249
transform -1 0 56544 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2233_
timestamp 1683973020
transform 1 0 55008 0 -1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _2234_
timestamp 1676557249
transform -1 0 59136 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2235_
timestamp 1683973020
transform 1 0 58176 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2236_
timestamp 1676557249
transform -1 0 61440 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2237_
timestamp 1683973020
transform 1 0 60288 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2238_
timestamp 1676557249
transform -1 0 61056 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2239_
timestamp 1683973020
transform 1 0 60096 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2240_
timestamp 1676557249
transform 1 0 60000 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2241_
timestamp 1683973020
transform -1 0 60096 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2242_
timestamp 1676557249
transform -1 0 56064 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2243_
timestamp 1683973020
transform 1 0 55296 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2244_
timestamp 1676557249
transform -1 0 57024 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2245_
timestamp 1683973020
transform 1 0 56160 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2246_
timestamp 1676557249
transform -1 0 56736 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2247_
timestamp 1683973020
transform 1 0 55872 0 -1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2248_
timestamp 1676557249
transform -1 0 55104 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2249_
timestamp 1683973020
transform -1 0 55584 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2250_
timestamp 1676557249
transform 1 0 51552 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2251_
timestamp 1683973020
transform -1 0 52416 0 -1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _2252_
timestamp 1676557249
transform -1 0 47424 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2253_
timestamp 1683973020
transform 1 0 45600 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2254_
timestamp 1676557249
transform 1 0 51168 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2255_
timestamp 1683973020
transform 1 0 51072 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2256_
timestamp 1676557249
transform -1 0 51456 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2257_
timestamp 1683973020
transform -1 0 51264 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2258_
timestamp 1676557249
transform -1 0 52320 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2259_
timestamp 1683973020
transform 1 0 51456 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2260_
timestamp 1676557249
transform -1 0 52800 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2261_
timestamp 1683973020
transform 1 0 52032 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2262_
timestamp 1676557249
transform -1 0 51840 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2263_
timestamp 1683973020
transform 1 0 50976 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2264_
timestamp 1676557249
transform -1 0 50496 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2265_
timestamp 1683973020
transform -1 0 51264 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2266_
timestamp 1676557249
transform 1 0 45504 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2267_
timestamp 1683973020
transform 1 0 45408 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _2268_
timestamp 1676557249
transform 1 0 45408 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2269_
timestamp 1683973020
transform -1 0 46272 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2270_
timestamp 1676557249
transform 1 0 46656 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2271_
timestamp 1683973020
transform 1 0 47040 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2272_
timestamp 1676557249
transform -1 0 47904 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2273_
timestamp 1683973020
transform 1 0 47040 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2274_
timestamp 1676557249
transform -1 0 46464 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _2275_
timestamp 1683973020
transform -1 0 46656 0 -1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2276_
timestamp 1676557249
transform 1 0 43200 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2277_
timestamp 1683973020
transform -1 0 44064 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2278_
timestamp 1676557249
transform 1 0 41472 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2279_
timestamp 1683973020
transform -1 0 42432 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2280_
timestamp 1676557249
transform -1 0 41664 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2281_
timestamp 1683973020
transform -1 0 41760 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2282_
timestamp 1676557249
transform -1 0 41184 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2283_
timestamp 1683973020
transform 1 0 40320 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2284_
timestamp 1676557249
transform -1 0 41376 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2285_
timestamp 1683973020
transform 1 0 40512 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2286_
timestamp 1676557249
transform -1 0 36960 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2287_
timestamp 1683973020
transform 1 0 36096 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2288_
timestamp 1676557249
transform 1 0 35232 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2289_
timestamp 1683973020
transform -1 0 35904 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2290_
timestamp 1676557249
transform -1 0 33504 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2291_
timestamp 1683973020
transform 1 0 32640 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2292_
timestamp 1676557249
transform 1 0 31968 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2293_
timestamp 1683973020
transform 1 0 31776 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2294_
timestamp 1676557249
transform 1 0 28800 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2295_
timestamp 1683973020
transform 1 0 28608 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _2296_
timestamp 1676557249
transform -1 0 9696 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2297_
timestamp 1683973020
transform 1 0 8736 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2298_
timestamp 1676557249
transform 1 0 4320 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2299_
timestamp 1683973020
transform -1 0 5184 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2300_
timestamp 1676557249
transform 1 0 3744 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2301_
timestamp 1683973020
transform -1 0 6432 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2302_
timestamp 1676557249
transform -1 0 5280 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2303_
timestamp 1683973020
transform 1 0 4512 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2304_
timestamp 1676557249
transform -1 0 5088 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2305_
timestamp 1683973020
transform -1 0 4704 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2306_
timestamp 1676557249
transform -1 0 5184 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2307_
timestamp 1683973020
transform 1 0 4416 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2308_
timestamp 1676557249
transform -1 0 5376 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2309_
timestamp 1683973020
transform 1 0 4416 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2310_
timestamp 1676557249
transform -1 0 4992 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2311_
timestamp 1683973020
transform -1 0 4608 0 -1 15876
box -48 -56 528 834
use sg13g2_tiehi  _2312__327
timestamp 1680000651
transform -1 0 23616 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2312_
timestamp 1746535128
transform 1 0 22752 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2313__326
timestamp 1680000651
transform 1 0 25632 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2313_
timestamp 1746535128
transform 1 0 26016 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2314__324
timestamp 1680000651
transform -1 0 30048 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2314_
timestamp 1746535128
transform 1 0 29184 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2315_
timestamp 1746535128
transform 1 0 32256 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2315__322
timestamp 1680000651
transform -1 0 33120 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  _2316__320
timestamp 1680000651
transform -1 0 36096 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2316_
timestamp 1746535128
transform 1 0 35328 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2317__318
timestamp 1680000651
transform -1 0 39840 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2317_
timestamp 1746535128
transform 1 0 38688 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2318__316
timestamp 1680000651
transform 1 0 41472 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2318_
timestamp 1746535128
transform 1 0 41376 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2319__314
timestamp 1680000651
transform -1 0 40608 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2319_
timestamp 1746535128
transform 1 0 39744 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2320_
timestamp 1746535128
transform 1 0 40224 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2320__312
timestamp 1680000651
transform -1 0 41088 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2321__310
timestamp 1680000651
transform 1 0 37920 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2321_
timestamp 1746535128
transform -1 0 39936 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2322_
timestamp 1746535128
transform -1 0 37440 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2322__308
timestamp 1680000651
transform 1 0 35328 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2323_
timestamp 1746535128
transform 1 0 30912 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2323__306
timestamp 1680000651
transform -1 0 31776 0 -1 15876
box -48 -56 432 834
use sg13g2_tiehi  _2324__304
timestamp 1680000651
transform -1 0 33792 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2324_
timestamp 1746535128
transform 1 0 32928 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2325_
timestamp 1746535128
transform 1 0 33792 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2325__302
timestamp 1680000651
transform -1 0 34656 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2326__300
timestamp 1680000651
transform 1 0 35904 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2326_
timestamp 1746535128
transform 1 0 36288 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2327__298
timestamp 1680000651
transform -1 0 40128 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2327_
timestamp 1746535128
transform 1 0 39264 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2328__296
timestamp 1680000651
transform 1 0 41184 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2328_
timestamp 1746535128
transform 1 0 41472 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2329__294
timestamp 1680000651
transform -1 0 45024 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2329_
timestamp 1746535128
transform 1 0 44160 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2330__292
timestamp 1680000651
transform -1 0 46176 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2330_
timestamp 1746535128
transform 1 0 45312 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2331__290
timestamp 1680000651
transform -1 0 46464 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2331_
timestamp 1746535128
transform 1 0 45600 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2332__288
timestamp 1680000651
transform -1 0 50400 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2332_
timestamp 1746535128
transform 1 0 49536 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2333__286
timestamp 1680000651
transform -1 0 52224 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2333_
timestamp 1746535128
transform 1 0 51360 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2334__284
timestamp 1680000651
transform -1 0 51264 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2334_
timestamp 1746535128
transform 1 0 50400 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2335_
timestamp 1746535128
transform 1 0 49824 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2335__282
timestamp 1680000651
transform 1 0 50112 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2336_
timestamp 1746535128
transform 1 0 48000 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2336__280
timestamp 1680000651
transform 1 0 47616 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2337_
timestamp 1746535128
transform 1 0 45408 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2337__278
timestamp 1680000651
transform -1 0 46272 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2338__276
timestamp 1680000651
transform -1 0 45408 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2338_
timestamp 1746535128
transform 1 0 44544 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2339__274
timestamp 1680000651
transform -1 0 44064 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2339_
timestamp 1746535128
transform 1 0 43200 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2340__272
timestamp 1680000651
transform -1 0 47136 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2340_
timestamp 1746535128
transform 1 0 46272 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2341__270
timestamp 1680000651
transform -1 0 49440 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2341_
timestamp 1746535128
transform 1 0 48576 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2342_
timestamp 1746535128
transform 1 0 50688 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2342__268
timestamp 1680000651
transform 1 0 50688 0 -1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2343__266
timestamp 1680000651
transform -1 0 54624 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2343_
timestamp 1746535128
transform 1 0 53760 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2344_
timestamp 1746535128
transform 1 0 54816 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2344__264
timestamp 1680000651
transform -1 0 55680 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2345__262
timestamp 1680000651
transform 1 0 56064 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2345_
timestamp 1746535128
transform 1 0 56352 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2346__260
timestamp 1680000651
transform -1 0 56736 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2346_
timestamp 1746535128
transform 1 0 55872 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2347_
timestamp 1746535128
transform 1 0 56736 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2347__258
timestamp 1680000651
transform -1 0 57600 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2348__256
timestamp 1680000651
transform -1 0 60000 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2348_
timestamp 1746535128
transform 1 0 58752 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2349__254
timestamp 1680000651
transform 1 0 54816 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2349_
timestamp 1746535128
transform -1 0 56256 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2350__252
timestamp 1680000651
transform -1 0 54240 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2350_
timestamp 1746535128
transform 1 0 53376 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2351__250
timestamp 1680000651
transform -1 0 61152 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2351_
timestamp 1746535128
transform 1 0 59136 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2352__248
timestamp 1680000651
transform -1 0 62496 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2352_
timestamp 1746535128
transform 1 0 61728 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2353_
timestamp 1746535128
transform 1 0 62784 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2353__246
timestamp 1680000651
transform -1 0 63648 0 -1 3780
box -48 -56 432 834
use sg13g2_tiehi  _2354__244
timestamp 1680000651
transform -1 0 63744 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2354_
timestamp 1746535128
transform 1 0 62880 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2355__242
timestamp 1680000651
transform -1 0 63360 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2355_
timestamp 1746535128
transform 1 0 62112 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2356__240
timestamp 1680000651
transform 1 0 62112 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2356_
timestamp 1746535128
transform 1 0 62112 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2357__238
timestamp 1680000651
transform 1 0 61824 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2357_
timestamp 1746535128
transform -1 0 63456 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2358_
timestamp 1746535128
transform 1 0 61152 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2358__236
timestamp 1680000651
transform -1 0 62784 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2359_
timestamp 1746535128
transform 1 0 64608 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2359__234
timestamp 1680000651
transform -1 0 65472 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2360__232
timestamp 1680000651
transform -1 0 68352 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2360_
timestamp 1746535128
transform 1 0 67488 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2361_
timestamp 1746535128
transform 1 0 67296 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2361__230
timestamp 1680000651
transform 1 0 67296 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2362__228
timestamp 1680000651
transform -1 0 68160 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2362_
timestamp 1746535128
transform 1 0 66816 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2363__226
timestamp 1680000651
transform 1 0 68256 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2363_
timestamp 1746535128
transform 1 0 68544 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2364__224
timestamp 1680000651
transform 1 0 69120 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2364_
timestamp 1746535128
transform 1 0 69120 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2365__222
timestamp 1680000651
transform -1 0 66816 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2365_
timestamp 1746535128
transform 1 0 65952 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2366__220
timestamp 1680000651
transform 1 0 69216 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2366_
timestamp 1746535128
transform 1 0 68928 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2367__218
timestamp 1680000651
transform 1 0 70656 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2367_
timestamp 1746535128
transform 1 0 71328 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2368__216
timestamp 1680000651
transform 1 0 75744 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2368_
timestamp 1746535128
transform 1 0 75552 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2369__214
timestamp 1680000651
transform 1 0 74208 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2369_
timestamp 1746535128
transform 1 0 74400 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2370__212
timestamp 1680000651
transform 1 0 74496 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2370_
timestamp 1746535128
transform -1 0 76128 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2371__210
timestamp 1680000651
transform -1 0 74592 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2371_
timestamp 1746535128
transform 1 0 73440 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2372_
timestamp 1746535128
transform 1 0 73344 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2372__208
timestamp 1680000651
transform -1 0 74208 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2373_
timestamp 1746535128
transform 1 0 72384 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2373__206
timestamp 1680000651
transform -1 0 73248 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2374__204
timestamp 1680000651
transform 1 0 71712 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2374_
timestamp 1746535128
transform 1 0 72096 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2375__202
timestamp 1680000651
transform -1 0 72960 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2375_
timestamp 1746535128
transform 1 0 72096 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2376__456
timestamp 1680000651
transform 1 0 73152 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2376_
timestamp 1746535128
transform 1 0 73152 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2377__454
timestamp 1680000651
transform -1 0 73824 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2377_
timestamp 1746535128
transform 1 0 72960 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2378__452
timestamp 1680000651
transform -1 0 74208 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2378_
timestamp 1746535128
transform 1 0 73344 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2379__450
timestamp 1680000651
transform -1 0 74400 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2379_
timestamp 1746535128
transform 1 0 73536 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2380__448
timestamp 1680000651
transform 1 0 74784 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2380_
timestamp 1746535128
transform 1 0 74688 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2381__446
timestamp 1680000651
transform -1 0 74976 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2381_
timestamp 1746535128
transform 1 0 74112 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2382__444
timestamp 1680000651
transform -1 0 76320 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2382_
timestamp 1746535128
transform 1 0 75456 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2383__442
timestamp 1680000651
transform 1 0 71712 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2383_
timestamp 1746535128
transform -1 0 73440 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2384__440
timestamp 1680000651
transform 1 0 69216 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2384_
timestamp 1746535128
transform -1 0 71424 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2385__438
timestamp 1680000651
transform -1 0 66528 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2385_
timestamp 1746535128
transform 1 0 65664 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2386_
timestamp 1746535128
transform 1 0 64128 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2386__436
timestamp 1680000651
transform -1 0 64992 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  _2387__434
timestamp 1680000651
transform -1 0 66912 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2387_
timestamp 1746535128
transform 1 0 66144 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2388__432
timestamp 1680000651
transform -1 0 70080 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2388_
timestamp 1746535128
transform 1 0 69216 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2389__430
timestamp 1680000651
transform -1 0 69120 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2389_
timestamp 1746535128
transform 1 0 68160 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2390__428
timestamp 1680000651
transform 1 0 67200 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2390_
timestamp 1746535128
transform 1 0 67584 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2391__426
timestamp 1680000651
transform 1 0 69120 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2391_
timestamp 1746535128
transform 1 0 69120 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2392_
timestamp 1746535128
transform -1 0 68160 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2392__424
timestamp 1680000651
transform 1 0 66144 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2393__422
timestamp 1680000651
transform -1 0 62400 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2393_
timestamp 1746535128
transform 1 0 61536 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2394__420
timestamp 1680000651
transform -1 0 62688 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2394_
timestamp 1746535128
transform 1 0 61824 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2395__418
timestamp 1680000651
transform -1 0 63936 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2395_
timestamp 1746535128
transform 1 0 63072 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2396__416
timestamp 1680000651
transform -1 0 61632 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2396_
timestamp 1746535128
transform 1 0 60288 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2397__414
timestamp 1680000651
transform -1 0 60576 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2397_
timestamp 1746535128
transform 1 0 59712 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2398__412
timestamp 1680000651
transform 1 0 61632 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2398_
timestamp 1746535128
transform 1 0 61632 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2399__410
timestamp 1680000651
transform -1 0 56736 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2399_
timestamp 1746535128
transform 1 0 55872 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2400__408
timestamp 1680000651
transform -1 0 55200 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2400_
timestamp 1746535128
transform 1 0 54336 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2401__406
timestamp 1680000651
transform -1 0 58944 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2401_
timestamp 1746535128
transform 1 0 57888 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2402_
timestamp 1746535128
transform 1 0 57696 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2402__404
timestamp 1680000651
transform -1 0 58560 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  _2403__402
timestamp 1680000651
transform -1 0 58080 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2403_
timestamp 1746535128
transform 1 0 57216 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2404__400
timestamp 1680000651
transform -1 0 58272 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2404_
timestamp 1746535128
transform 1 0 57408 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2405__398
timestamp 1680000651
transform -1 0 56448 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2405_
timestamp 1746535128
transform -1 0 56736 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2406_
timestamp 1746535128
transform 1 0 52800 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2406__396
timestamp 1680000651
transform 1 0 52032 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2407_
timestamp 1746535128
transform 1 0 52704 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2407__394
timestamp 1680000651
transform -1 0 53568 0 -1 30996
box -48 -56 432 834
use sg13g2_tiehi  _2408__392
timestamp 1680000651
transform -1 0 52992 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2408_
timestamp 1746535128
transform 1 0 52128 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2409__390
timestamp 1680000651
transform 1 0 48864 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2409_
timestamp 1746535128
transform -1 0 50976 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2410__388
timestamp 1680000651
transform 1 0 45696 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2410_
timestamp 1746535128
transform 1 0 46080 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2411__386
timestamp 1680000651
transform 1 0 47808 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2411_
timestamp 1746535128
transform 1 0 48192 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2412_
timestamp 1746535128
transform 1 0 48000 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2412__384
timestamp 1680000651
transform 1 0 48096 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  _2413__382
timestamp 1680000651
transform -1 0 49632 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2413_
timestamp 1746535128
transform 1 0 48768 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2414__380
timestamp 1680000651
transform 1 0 47136 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2414_
timestamp 1746535128
transform 1 0 48768 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2415__378
timestamp 1680000651
transform -1 0 48768 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2415_
timestamp 1746535128
transform 1 0 47904 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2416__376
timestamp 1680000651
transform -1 0 48480 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2416_
timestamp 1746535128
transform 1 0 47616 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2417__374
timestamp 1680000651
transform -1 0 43104 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2417_
timestamp 1746535128
transform 1 0 42240 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2418__372
timestamp 1680000651
transform -1 0 43104 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2418_
timestamp 1746535128
transform 1 0 42240 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2419_
timestamp 1746535128
transform 1 0 43776 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2419__370
timestamp 1680000651
transform 1 0 43584 0 1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2420__368
timestamp 1680000651
transform 1 0 44448 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2420_
timestamp 1746535128
transform -1 0 46080 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2421__366
timestamp 1680000651
transform -1 0 44736 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2421_
timestamp 1746535128
transform 1 0 43488 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2422__364
timestamp 1680000651
transform -1 0 40896 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2422_
timestamp 1746535128
transform 1 0 40032 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2423__362
timestamp 1680000651
transform -1 0 39264 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2423_
timestamp 1746535128
transform 1 0 38400 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2424_
timestamp 1746535128
transform 1 0 37728 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2424__360
timestamp 1680000651
transform -1 0 38592 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2425_
timestamp 1746535128
transform 1 0 37152 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2425__358
timestamp 1680000651
transform -1 0 38016 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2426_
timestamp 1746535128
transform 1 0 38400 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2426__356
timestamp 1680000651
transform 1 0 38592 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2427_
timestamp 1746535128
transform 1 0 35040 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2427__354
timestamp 1680000651
transform 1 0 35232 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2428_
timestamp 1746535128
transform -1 0 34464 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2428__352
timestamp 1680000651
transform 1 0 32448 0 1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2429__350
timestamp 1680000651
transform -1 0 30624 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2429_
timestamp 1746535128
transform 1 0 29760 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2430__348
timestamp 1680000651
transform -1 0 28992 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2430_
timestamp 1746535128
transform 1 0 28128 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2431_
timestamp 1746535128
transform -1 0 28320 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2431__346
timestamp 1680000651
transform 1 0 26208 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  _2432__344
timestamp 1680000651
transform 1 0 6336 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2432_
timestamp 1746535128
transform -1 0 8448 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2433__342
timestamp 1680000651
transform -1 0 2112 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2433_
timestamp 1746535128
transform 1 0 1248 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2434__340
timestamp 1680000651
transform -1 0 2016 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2434_
timestamp 1746535128
transform 1 0 1152 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2435__338
timestamp 1680000651
transform 1 0 1344 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2435_
timestamp 1746535128
transform 1 0 1440 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2436__336
timestamp 1680000651
transform 1 0 1056 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2436_
timestamp 1746535128
transform 1 0 1056 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2437_
timestamp 1746535128
transform 1 0 1440 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2437__334
timestamp 1680000651
transform 1 0 1536 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2438_
timestamp 1746535128
transform 1 0 2016 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2438__332
timestamp 1680000651
transform -1 0 3168 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2439_
timestamp 1746535128
transform 1 0 960 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2439__330
timestamp 1680000651
transform -1 0 1824 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2440_
timestamp 1746535128
transform 1 0 23040 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2440__328
timestamp 1680000651
transform -1 0 24000 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2441__325
timestamp 1680000651
transform -1 0 28032 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2441_
timestamp 1746535128
transform 1 0 27168 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2442_
timestamp 1746535128
transform 1 0 30336 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2442__321
timestamp 1680000651
transform -1 0 31200 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2443__317
timestamp 1680000651
transform -1 0 34176 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2443_
timestamp 1746535128
transform 1 0 32928 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2444_
timestamp 1746535128
transform 1 0 36096 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2444__313
timestamp 1680000651
transform -1 0 37056 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2445__309
timestamp 1680000651
transform -1 0 40992 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2445_
timestamp 1746535128
transform 1 0 38688 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2446__305
timestamp 1680000651
transform -1 0 45024 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2446_
timestamp 1746535128
transform 1 0 43680 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2447_
timestamp 1746535128
transform 1 0 43104 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2447__301
timestamp 1680000651
transform -1 0 43968 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2448__297
timestamp 1680000651
transform -1 0 44160 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2448_
timestamp 1746535128
transform 1 0 43008 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2449__293
timestamp 1680000651
transform -1 0 41184 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2449_
timestamp 1746535128
transform 1 0 40224 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2450__289
timestamp 1680000651
transform -1 0 38112 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2450_
timestamp 1746535128
transform 1 0 37248 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2451__285
timestamp 1680000651
transform -1 0 35040 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2451_
timestamp 1746535128
transform 1 0 34176 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2452_
timestamp 1746535128
transform 1 0 29856 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2452__281
timestamp 1680000651
transform -1 0 30720 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2453_
timestamp 1746535128
transform 1 0 36864 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2453__277
timestamp 1680000651
transform -1 0 37728 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2454__273
timestamp 1680000651
transform -1 0 39840 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2454_
timestamp 1746535128
transform 1 0 38976 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2455__269
timestamp 1680000651
transform -1 0 43104 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2455_
timestamp 1746535128
transform 1 0 42240 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2456__265
timestamp 1680000651
transform -1 0 45216 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2456_
timestamp 1746535128
transform 1 0 44064 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2457_
timestamp 1746535128
transform 1 0 46656 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2457__261
timestamp 1680000651
transform -1 0 47520 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2458__257
timestamp 1680000651
transform -1 0 49632 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2458_
timestamp 1746535128
transform 1 0 48672 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2459__253
timestamp 1680000651
transform -1 0 49728 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2459_
timestamp 1746535128
transform 1 0 48768 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2460__249
timestamp 1680000651
transform -1 0 53184 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2460_
timestamp 1746535128
transform 1 0 52224 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2461__245
timestamp 1680000651
transform -1 0 55392 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2461_
timestamp 1746535128
transform 1 0 54528 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2462__241
timestamp 1680000651
transform -1 0 55200 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2462_
timestamp 1746535128
transform 1 0 54336 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2463_
timestamp 1746535128
transform 1 0 53760 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2463__237
timestamp 1680000651
transform -1 0 54624 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2464_
timestamp 1746535128
transform 1 0 51936 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2464__233
timestamp 1680000651
transform -1 0 52800 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2465_
timestamp 1746535128
transform 1 0 49344 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2465__229
timestamp 1680000651
transform -1 0 50208 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2466__225
timestamp 1680000651
transform -1 0 48768 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2466_
timestamp 1746535128
transform 1 0 47904 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2467_
timestamp 1746535128
transform 1 0 46176 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2467__221
timestamp 1680000651
transform -1 0 47136 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  _2468__217
timestamp 1680000651
transform -1 0 50400 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2468_
timestamp 1746535128
transform 1 0 49536 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2469__213
timestamp 1680000651
transform -1 0 51072 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2469_
timestamp 1746535128
transform 1 0 50208 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2470_
timestamp 1746535128
transform 1 0 53088 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2470__209
timestamp 1680000651
transform -1 0 53952 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  _2471__205
timestamp 1680000651
transform -1 0 57888 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2471_
timestamp 1746535128
transform 1 0 57024 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2472__201
timestamp 1680000651
transform -1 0 58944 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2472_
timestamp 1746535128
transform 1 0 58080 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2473__453
timestamp 1680000651
transform -1 0 60096 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2473_
timestamp 1746535128
transform 1 0 59232 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2474__449
timestamp 1680000651
transform -1 0 60576 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2474_
timestamp 1746535128
transform 1 0 59520 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2475__445
timestamp 1680000651
transform -1 0 61248 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2475_
timestamp 1746535128
transform 1 0 60384 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2476_
timestamp 1746535128
transform 1 0 61152 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2476__441
timestamp 1680000651
transform -1 0 62016 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2477__437
timestamp 1680000651
transform -1 0 56928 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2477_
timestamp 1746535128
transform 1 0 56064 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2478__433
timestamp 1680000651
transform -1 0 57696 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2478_
timestamp 1746535128
transform 1 0 56544 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2479__429
timestamp 1680000651
transform -1 0 60480 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2479_
timestamp 1746535128
transform 1 0 59616 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2480__425
timestamp 1680000651
transform -1 0 65376 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2480_
timestamp 1746535128
transform 1 0 64416 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2481__421
timestamp 1680000651
transform -1 0 67200 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2481_
timestamp 1746535128
transform 1 0 66336 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2482__417
timestamp 1680000651
transform -1 0 67488 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2482_
timestamp 1746535128
transform 1 0 66528 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2483__413
timestamp 1680000651
transform -1 0 66816 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2483_
timestamp 1746535128
transform 1 0 65952 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2484__409
timestamp 1680000651
transform -1 0 66144 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2484_
timestamp 1746535128
transform 1 0 65184 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2485_
timestamp 1746535128
transform 1 0 64704 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2485__405
timestamp 1680000651
transform -1 0 65664 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2486_
timestamp 1746535128
transform 1 0 60480 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2486__401
timestamp 1680000651
transform -1 0 61344 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2487_
timestamp 1746535128
transform 1 0 65376 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2487__397
timestamp 1680000651
transform -1 0 66240 0 1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2488__393
timestamp 1680000651
transform -1 0 71616 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2488_
timestamp 1746535128
transform 1 0 70272 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2489__389
timestamp 1680000651
transform -1 0 71328 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2489_
timestamp 1746535128
transform 1 0 70368 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2490__385
timestamp 1680000651
transform -1 0 71616 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2490_
timestamp 1746535128
transform 1 0 70368 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2491__381
timestamp 1680000651
transform -1 0 72480 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2491_
timestamp 1746535128
transform 1 0 71616 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2492__377
timestamp 1680000651
transform -1 0 72768 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2492_
timestamp 1746535128
transform 1 0 71904 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2493__373
timestamp 1680000651
transform -1 0 69696 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2493_
timestamp 1746535128
transform 1 0 68736 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2494__369
timestamp 1680000651
transform -1 0 72672 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2494_
timestamp 1746535128
transform 1 0 71808 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2495__365
timestamp 1680000651
transform -1 0 74976 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2495_
timestamp 1746535128
transform 1 0 73152 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2496__361
timestamp 1680000651
transform 1 0 77952 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2496_
timestamp 1746535128
transform -1 0 79584 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2497__357
timestamp 1680000651
transform -1 0 78144 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2497_
timestamp 1746535128
transform 1 0 76992 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2498__353
timestamp 1680000651
transform -1 0 78144 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2498_
timestamp 1746535128
transform 1 0 76992 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2499_
timestamp 1746535128
transform 1 0 76992 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2499__349
timestamp 1680000651
transform -1 0 78048 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2500__345
timestamp 1680000651
transform -1 0 77952 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2500_
timestamp 1746535128
transform 1 0 76992 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2501_
timestamp 1746535128
transform 1 0 76800 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2501__341
timestamp 1680000651
transform -1 0 77664 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2502_
timestamp 1746535128
transform 1 0 76896 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2502__337
timestamp 1680000651
transform -1 0 77760 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2503__333
timestamp 1680000651
transform -1 0 76992 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2503_
timestamp 1746535128
transform 1 0 76128 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2504_
timestamp 1746535128
transform 1 0 76608 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2504__329
timestamp 1680000651
transform -1 0 77472 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2505__323
timestamp 1680000651
transform -1 0 77856 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2505_
timestamp 1746535128
transform 1 0 76992 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2506__315
timestamp 1680000651
transform -1 0 77856 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2506_
timestamp 1746535128
transform 1 0 76992 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2507_
timestamp 1746535128
transform 1 0 76992 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2507__307
timestamp 1680000651
transform -1 0 78144 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  _2508__299
timestamp 1680000651
transform -1 0 78144 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2508_
timestamp 1746535128
transform 1 0 76992 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2509__291
timestamp 1680000651
transform -1 0 78144 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2509_
timestamp 1746535128
transform 1 0 76992 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2510__283
timestamp 1680000651
transform -1 0 78816 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2510_
timestamp 1746535128
transform 1 0 76992 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2511__275
timestamp 1680000651
transform -1 0 74304 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2511_
timestamp 1746535128
transform 1 0 73440 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2512__267
timestamp 1680000651
transform -1 0 73056 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2512_
timestamp 1746535128
transform 1 0 72096 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2513_
timestamp 1746535128
transform 1 0 69024 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2513__259
timestamp 1680000651
transform -1 0 69984 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2514_
timestamp 1746535128
transform 1 0 67392 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2514__251
timestamp 1680000651
transform -1 0 68256 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2515_
timestamp 1746535128
transform 1 0 66624 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2515__243
timestamp 1680000651
transform -1 0 67584 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2516_
timestamp 1746535128
transform 1 0 72096 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2516__235
timestamp 1680000651
transform -1 0 73152 0 -1 32508
box -48 -56 432 834
use sg13g2_tiehi  _2517__227
timestamp 1680000651
transform -1 0 72576 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2517_
timestamp 1746535128
transform 1 0 71712 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2518_
timestamp 1746535128
transform 1 0 71328 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2518__219
timestamp 1680000651
transform -1 0 72192 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2519_
timestamp 1746535128
transform 1 0 70560 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2519__211
timestamp 1680000651
transform -1 0 71520 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2520_
timestamp 1746535128
transform 1 0 67872 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2520__203
timestamp 1680000651
transform -1 0 68832 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2521_
timestamp 1746535128
transform 1 0 63936 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2521__451
timestamp 1680000651
transform -1 0 65088 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2522_
timestamp 1746535128
transform 1 0 65664 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2522__443
timestamp 1680000651
transform -1 0 66528 0 -1 27972
box -48 -56 432 834
use sg13g2_tiehi  _2523__435
timestamp 1680000651
transform -1 0 66816 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2523_
timestamp 1746535128
transform 1 0 65952 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2524__427
timestamp 1680000651
transform -1 0 64032 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2524_
timestamp 1746535128
transform 1 0 63168 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2525__419
timestamp 1680000651
transform -1 0 63840 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2525_
timestamp 1746535128
transform 1 0 62976 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2526__411
timestamp 1680000651
transform 1 0 64320 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2526_
timestamp 1746535128
transform 1 0 64224 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2527__403
timestamp 1680000651
transform -1 0 60480 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2527_
timestamp 1746535128
transform 1 0 59040 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2528_
timestamp 1746535128
transform 1 0 55488 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2528__395
timestamp 1680000651
transform -1 0 56832 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  _2529__387
timestamp 1680000651
transform -1 0 59520 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2529_
timestamp 1746535128
transform 1 0 58656 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2530__379
timestamp 1680000651
transform -1 0 61440 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2530_
timestamp 1746535128
transform 1 0 60576 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2531_
timestamp 1746535128
transform 1 0 60480 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2531__371
timestamp 1680000651
transform -1 0 61440 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2532_
timestamp 1746535128
transform 1 0 60096 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2532__363
timestamp 1680000651
transform -1 0 61152 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2533__355
timestamp 1680000651
transform 1 0 55296 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2533_
timestamp 1746535128
transform 1 0 55008 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2534__347
timestamp 1680000651
transform -1 0 56928 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2534_
timestamp 1746535128
transform 1 0 56064 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2535__339
timestamp 1680000651
transform -1 0 56928 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2535_
timestamp 1746535128
transform 1 0 56064 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2536__331
timestamp 1680000651
transform -1 0 56448 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2536_
timestamp 1746535128
transform 1 0 55584 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2537_
timestamp 1746535128
transform 1 0 51936 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2537__319
timestamp 1680000651
transform -1 0 52800 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  _2538__303
timestamp 1680000651
transform 1 0 45984 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2538_
timestamp 1746535128
transform 1 0 45792 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2539__287
timestamp 1680000651
transform -1 0 51936 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2539_
timestamp 1746535128
transform 1 0 51072 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2540__271
timestamp 1680000651
transform -1 0 52608 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2540_
timestamp 1746535128
transform 1 0 51168 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2541__255
timestamp 1680000651
transform -1 0 52800 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2541_
timestamp 1746535128
transform 1 0 51936 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2542__239
timestamp 1680000651
transform -1 0 53184 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2542_
timestamp 1746535128
transform 1 0 52320 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2543__223
timestamp 1680000651
transform -1 0 52896 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2543_
timestamp 1746535128
transform 1 0 51648 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2544__207
timestamp 1680000651
transform -1 0 51648 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2544_
timestamp 1746535128
transform 1 0 50208 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2545__447
timestamp 1680000651
transform -1 0 46752 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2545_
timestamp 1746535128
transform 1 0 45888 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2546__431
timestamp 1680000651
transform -1 0 47232 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2546_
timestamp 1746535128
transform 1 0 46368 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2547_
timestamp 1746535128
transform 1 0 47040 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2547__415
timestamp 1680000651
transform -1 0 47904 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2548__399
timestamp 1680000651
transform -1 0 47904 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2548_
timestamp 1746535128
transform 1 0 47040 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2549__383
timestamp 1680000651
transform -1 0 47328 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2549_
timestamp 1746535128
transform 1 0 46464 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2550__367
timestamp 1680000651
transform -1 0 44256 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2550_
timestamp 1746535128
transform 1 0 43200 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2551__351
timestamp 1680000651
transform -1 0 42816 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2551_
timestamp 1746535128
transform 1 0 41856 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2552_
timestamp 1746535128
transform 1 0 41664 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2552__335
timestamp 1680000651
transform -1 0 42528 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2553__311
timestamp 1680000651
transform -1 0 41664 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2553_
timestamp 1746535128
transform 1 0 40800 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2554__279
timestamp 1680000651
transform -1 0 42336 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2554_
timestamp 1746535128
transform 1 0 40992 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2555_
timestamp 1746535128
transform 1 0 35712 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2555__247
timestamp 1680000651
transform 1 0 35328 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2556_
timestamp 1746535128
transform 1 0 35616 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2556__215
timestamp 1680000651
transform -1 0 36576 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2557_
timestamp 1746535128
transform 1 0 33024 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2557__439
timestamp 1680000651
transform -1 0 33888 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2558_
timestamp 1746535128
transform 1 0 32448 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2558__407
timestamp 1680000651
transform -1 0 33504 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2559_
timestamp 1746535128
transform 1 0 29184 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2559__375
timestamp 1680000651
transform -1 0 30144 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2560_
timestamp 1746535128
transform 1 0 9216 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2560__343
timestamp 1680000651
transform -1 0 10080 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  _2561__295
timestamp 1680000651
transform -1 0 6240 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2561_
timestamp 1746535128
transform 1 0 5184 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2562_
timestamp 1746535128
transform 1 0 4992 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2562__231
timestamp 1680000651
transform -1 0 5856 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2563_
timestamp 1746535128
transform 1 0 4992 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2563__423
timestamp 1680000651
transform -1 0 5856 0 1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2564__359
timestamp 1680000651
transform -1 0 5568 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2564_
timestamp 1746535128
transform 1 0 4704 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2565__263
timestamp 1680000651
transform -1 0 6240 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2565_
timestamp 1746535128
transform 1 0 4896 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2566_
timestamp 1746535128
transform 1 0 4992 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2566__391
timestamp 1680000651
transform -1 0 6528 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2567_
timestamp 1746535128
transform 1 0 4512 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2567__455
timestamp 1680000651
transform -1 0 5376 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2832_
timestamp 1676381911
transform -1 0 1824 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _2833_
timestamp 1676381911
transform -1 0 1824 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _2834_
timestamp 1676381911
transform -1 0 1440 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _2835_
timestamp 1676381911
transform -1 0 1536 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _2836_
timestamp 1676381911
transform -1 0 1440 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2837_
timestamp 1676381911
transform -1 0 1536 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2838_
timestamp 1676381911
transform -1 0 1440 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _2839_
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2840_
timestamp 1676381911
transform -1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _2841_
timestamp 1676381911
transform -1 0 1248 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _2842_
timestamp 1676381911
transform -1 0 1536 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _2843_
timestamp 1676381911
transform -1 0 1152 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _2844_
timestamp 1676381911
transform -1 0 1344 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _2845_
timestamp 1676381911
transform -1 0 1824 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _2846_
timestamp 1676381911
transform -1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2847_
timestamp 1676381911
transform -1 0 1824 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform -1 0 40704 0 -1 20412
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_0__f_clk
timestamp 1676553496
transform -1 0 52896 0 -1 9828
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_1__f_clk
timestamp 1676553496
transform 1 0 37248 0 -1 11340
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_2__f_clk
timestamp 1676553496
transform -1 0 55200 0 1 27972
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_3__f_clk
timestamp 1676553496
transform 1 0 44640 0 1 26460
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_leaf_0_clk
timestamp 1676451365
transform 1 0 4896 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_1_clk
timestamp 1676451365
transform -1 0 32352 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_2_clk
timestamp 1676451365
transform -1 0 37536 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_3_clk
timestamp 1676451365
transform 1 0 47520 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_4_clk
timestamp 1676451365
transform 1 0 49152 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_5_clk
timestamp 1676451365
transform -1 0 59712 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_6_clk
timestamp 1676451365
transform -1 0 71712 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_7_clk
timestamp 1676451365
transform 1 0 72576 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_8_clk
timestamp 1676451365
transform -1 0 70464 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_9_clk
timestamp 1676451365
transform -1 0 51744 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_10_clk
timestamp 1676451365
transform -1 0 52800 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_11_clk
timestamp 1676451365
transform 1 0 72000 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_12_clk
timestamp 1676451365
transform 1 0 71040 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_13_clk
timestamp 1676451365
transform -1 0 71040 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_14_clk
timestamp 1676451365
transform -1 0 60288 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_15_clk
timestamp 1676451365
transform -1 0 50400 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_16_clk
timestamp 1676451365
transform 1 0 45984 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_17_clk
timestamp 1676451365
transform 1 0 36960 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_18_clk
timestamp 1676451365
transform -1 0 5376 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkload0
timestamp 1676451365
transform -1 0 46176 0 1 24948
box -48 -56 1296 834
use sg13g2_inv_2  clkload1
timestamp 1676382947
transform 1 0 51552 0 1 15876
box -48 -56 432 834
use sg13g2_inv_2  clkload2
timestamp 1676382947
transform 1 0 72384 0 -1 3780
box -48 -56 432 834
use sg13g2_inv_2  clkload3
timestamp 1676382947
transform 1 0 48768 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_8  clkload4
timestamp 1676383150
transform 1 0 4896 0 -1 12852
box -48 -56 1008 834
use sg13g2_buf_8  clkload5
timestamp 1676451365
transform 1 0 45984 0 1 14364
box -48 -56 1296 834
use sg13g2_inv_8  clkload6
timestamp 1676383150
transform 1 0 36384 0 1 14364
box -48 -56 1008 834
use sg13g2_inv_16  clkload7
timestamp 1676383183
transform 1 0 4128 0 1 5292
box -48 -56 1872 834
use sg13g2_inv_1  clkload8
timestamp 1676382929
transform 1 0 36288 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  clkload9
timestamp 1676382929
transform -1 0 67584 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_4  clkload10
timestamp 1676383058
transform -1 0 72864 0 1 756
box -48 -56 624 834
use sg13g2_inv_1  clkload11
timestamp 1676382929
transform 1 0 47904 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  clkload12
timestamp 1676382929
transform 1 0 48384 0 -1 32508
box -48 -56 336 834
use dac128module  dac
timestamp 0
transform 1 0 53240 0 1 17400
box 0 0 1 1
use sg13g2_inv_1  digitalen.g\[0\].u.inv1
timestamp 1676382929
transform 1 0 52512 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[0\].u.inv2
timestamp 1676382929
transform -1 0 52800 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv1
timestamp 1676382929
transform 1 0 78816 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv2
timestamp 1676382929
transform 1 0 79296 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv1
timestamp 1676382929
transform 1 0 79008 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv2
timestamp 1676382929
transform 1 0 79296 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv1
timestamp 1676382929
transform 1 0 52512 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv2
timestamp 1676382929
transform -1 0 52224 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform 1 0 21504 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform 1 0 27936 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 2688 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform -1 0 41184 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform -1 0 47616 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform 1 0 49824 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform 1 0 43008 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform 1 0 38976 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform -1 0 41280 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 49920 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform 1 0 49248 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform 1 0 38784 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 57312 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform -1 0 57600 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform -1 0 68928 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 68640 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 60672 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform 1 0 58752 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform -1 0 71040 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform -1 0 67680 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 58272 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform 1 0 1920 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform -1 0 25728 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform 1 0 26208 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout47
timestamp 1676381911
transform 1 0 26784 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform -1 0 2976 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 41376 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout50
timestamp 1676381911
transform 1 0 49536 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform 1 0 48192 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout52
timestamp 1676381911
transform -1 0 42144 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform 1 0 39456 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 49248 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform 1 0 49344 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform 1 0 39072 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform 1 0 57312 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform -1 0 59040 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout59
timestamp 1676381911
transform -1 0 70368 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout60
timestamp 1676381911
transform 1 0 67104 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout61
timestamp 1676381911
transform 1 0 57888 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout62
timestamp 1676381911
transform 1 0 69408 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout63
timestamp 1676381911
transform -1 0 69120 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout64
timestamp 1676381911
transform -1 0 59040 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout65
timestamp 1676381911
transform 1 0 59520 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout66
timestamp 1676381911
transform 1 0 3168 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout67
timestamp 1676381911
transform 1 0 21408 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout68
timestamp 1676381911
transform 1 0 33312 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform -1 0 22176 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 9312 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform -1 0 45792 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform 1 0 44832 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform -1 0 50688 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform 1 0 44064 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform 1 0 40128 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform 1 0 51840 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform 1 0 48960 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform 1 0 42336 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 58656 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform -1 0 61728 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform -1 0 70272 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform -1 0 70848 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 60480 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform -1 0 60768 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform 1 0 71424 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 70368 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 60864 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform 1 0 8928 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform -1 0 3456 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform -1 0 4512 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform -1 0 32160 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout92
timestamp 1676381911
transform -1 0 37344 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout93
timestamp 1676381911
transform 1 0 24288 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout94
timestamp 1676381911
transform 1 0 31392 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout95
timestamp 1676381911
transform 1 0 36576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout96
timestamp 1676381911
transform 1 0 27072 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout97
timestamp 1676381911
transform -1 0 3840 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout98
timestamp 1676381911
transform 1 0 42048 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout99
timestamp 1676381911
transform 1 0 46464 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform -1 0 41760 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout101
timestamp 1676381911
transform -1 0 43200 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout102
timestamp 1676381911
transform 1 0 54624 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout103
timestamp 1676381911
transform -1 0 52032 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform -1 0 51456 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform 1 0 42816 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout106
timestamp 1676381911
transform 1 0 39456 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform -1 0 46368 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout108
timestamp 1676381911
transform 1 0 40320 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform -1 0 50496 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout110
timestamp 1676381911
transform 1 0 56160 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout111
timestamp 1676381911
transform -1 0 50112 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout112
timestamp 1676381911
transform 1 0 51072 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout113
timestamp 1676381911
transform 1 0 39936 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout114
timestamp 1676381911
transform 1 0 64704 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout115
timestamp 1676381911
transform -1 0 60192 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout116
timestamp 1676381911
transform -1 0 62112 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout117
timestamp 1676381911
transform -1 0 71232 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout118
timestamp 1676381911
transform 1 0 76416 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout119
timestamp 1676381911
transform 1 0 76416 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout120
timestamp 1676381911
transform 1 0 70464 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout121
timestamp 1676381911
transform -1 0 71232 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout122
timestamp 1676381911
transform 1 0 61632 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout123
timestamp 1676381911
transform 1 0 59136 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout124
timestamp 1676381911
transform -1 0 60672 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout125
timestamp 1676381911
transform -1 0 61344 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout126
timestamp 1676381911
transform -1 0 68928 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout127
timestamp 1676381911
transform -1 0 69408 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout128
timestamp 1676381911
transform -1 0 75168 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout129
timestamp 1676381911
transform 1 0 70848 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout130
timestamp 1676381911
transform 1 0 61344 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout131
timestamp 1676381911
transform 1 0 40512 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout132
timestamp 1676381911
transform 1 0 22176 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout133
timestamp 1676381911
transform 1 0 22176 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout134
timestamp 1676381911
transform -1 0 2688 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout135
timestamp 1676381911
transform 1 0 21888 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout136
timestamp 1676381911
transform -1 0 43584 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout137
timestamp 1676381911
transform 1 0 44448 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout138
timestamp 1676381911
transform 1 0 49824 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout139
timestamp 1676381911
transform 1 0 43584 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout140
timestamp 1676381911
transform -1 0 41088 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout141
timestamp 1676381911
transform 1 0 51840 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout142
timestamp 1676381911
transform 1 0 51456 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout143
timestamp 1676381911
transform -1 0 41760 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout144
timestamp 1676381911
transform -1 0 59520 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout145
timestamp 1676381911
transform -1 0 60864 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout146
timestamp 1676381911
transform -1 0 69792 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout147
timestamp 1676381911
transform -1 0 69984 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout148
timestamp 1676381911
transform 1 0 58656 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout149
timestamp 1676381911
transform -1 0 59136 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout150
timestamp 1676381911
transform 1 0 71040 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout151
timestamp 1676381911
transform 1 0 71712 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout152
timestamp 1676381911
transform 1 0 60480 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout153
timestamp 1676381911
transform 1 0 2688 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout154
timestamp 1676381911
transform -1 0 3936 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout155
timestamp 1676381911
transform 1 0 23904 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout156
timestamp 1676381911
transform 1 0 23520 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout157
timestamp 1676381911
transform -1 0 1920 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout158
timestamp 1676381911
transform -1 0 45408 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout159
timestamp 1676381911
transform -1 0 46752 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout160
timestamp 1676381911
transform -1 0 49440 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout161
timestamp 1676381911
transform 1 0 51552 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout162
timestamp 1676381911
transform 1 0 44256 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout163
timestamp 1676381911
transform 1 0 40608 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout164
timestamp 1676381911
transform 1 0 42048 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout165
timestamp 1676381911
transform -1 0 51456 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout166
timestamp 1676381911
transform 1 0 51552 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout167
timestamp 1676381911
transform 1 0 40320 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout168
timestamp 1676381911
transform 1 0 59424 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout169
timestamp 1676381911
transform -1 0 62880 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout170
timestamp 1676381911
transform 1 0 70272 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout171
timestamp 1676381911
transform -1 0 70848 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout172
timestamp 1676381911
transform 1 0 61440 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout173
timestamp 1676381911
transform -1 0 60768 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout174
timestamp 1676381911
transform -1 0 72192 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout175
timestamp 1676381911
transform -1 0 72480 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout176
timestamp 1676381911
transform 1 0 60288 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout177
timestamp 1676381911
transform 1 0 1920 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout178
timestamp 1676381911
transform -1 0 2784 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout179
timestamp 1676381911
transform 1 0 22272 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout180
timestamp 1676381911
transform 1 0 27360 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout181
timestamp 1676381911
transform -1 0 5856 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout182
timestamp 1676381911
transform -1 0 41568 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout183
timestamp 1676381911
transform -1 0 48000 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout184
timestamp 1676381911
transform 1 0 49344 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout185
timestamp 1676381911
transform -1 0 41856 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout186
timestamp 1676381911
transform -1 0 40224 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout187
timestamp 1676381911
transform 1 0 42336 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout188
timestamp 1676381911
transform -1 0 56928 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout189
timestamp 1676381911
transform -1 0 51072 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout190
timestamp 1676381911
transform 1 0 42720 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout191
timestamp 1676381911
transform 1 0 58176 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout192
timestamp 1676381911
transform 1 0 57792 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout193
timestamp 1676381911
transform 1 0 69408 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout194
timestamp 1676381911
transform -1 0 69312 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout195
timestamp 1676381911
transform 1 0 57216 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout196
timestamp 1676381911
transform -1 0 60096 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout197
timestamp 1676381911
transform 1 0 67488 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout198
timestamp 1676381911
transform -1 0 67968 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout199
timestamp 1676381911
transform 1 0 57600 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout200
timestamp 1676381911
transform 1 0 5856 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_567
timestamp 1679577901
transform 1 0 55008 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_576
timestamp 1677579658
transform 1 0 55872 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_602
timestamp 1677580104
transform 1 0 58368 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_631
timestamp 1679577901
transform 1 0 61152 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_635
timestamp 1677579658
transform 1 0 61536 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_651
timestamp 1679577901
transform 1 0 63072 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_655
timestamp 1677580104
transform 1 0 63456 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_675
timestamp 1679577901
transform 1 0 65376 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_679
timestamp 1677580104
transform 1 0 65760 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_713
timestamp 1677580104
transform 1 0 69024 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_715
timestamp 1677579658
transform 1 0 69216 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_720
timestamp 1677579658
transform 1 0 69696 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_753
timestamp 1677580104
transform 1 0 72864 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_755
timestamp 1677579658
transform 1 0 73056 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_783
timestamp 1677579658
transform 1 0 75744 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_789
timestamp 1679581782
transform 1 0 76320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_546
timestamp 1679577901
transform 1 0 52992 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_582
timestamp 1677579658
transform 1 0 56448 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_664
timestamp 1677579658
transform 1 0 64320 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_692
timestamp 1677580104
transform 1 0 67008 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_694
timestamp 1677579658
transform 1 0 67200 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_769
timestamp 1677579658
transform 1 0 74400 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_775
timestamp 1677579658
transform 1 0 74976 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_817
timestamp 1679577901
transform 1 0 79008 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_821
timestamp 1677580104
transform 1 0 79392 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_8
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_13
timestamp 1679577901
transform 1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_17
timestamp 1677580104
transform 1 0 2208 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_24
timestamp 1677579658
transform 1 0 2880 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_30
timestamp 1679581782
transform 1 0 3456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_37
timestamp 1679581782
transform 1 0 4128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_44
timestamp 1679581782
transform 1 0 4800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_51
timestamp 1679581782
transform 1 0 5472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_58
timestamp 1679581782
transform 1 0 6144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_65
timestamp 1679581782
transform 1 0 6816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_72
timestamp 1679581782
transform 1 0 7488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_79
timestamp 1679581782
transform 1 0 8160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_86
timestamp 1679581782
transform 1 0 8832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_93
timestamp 1679581782
transform 1 0 9504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_100
timestamp 1679581782
transform 1 0 10176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_107
timestamp 1679581782
transform 1 0 10848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_114
timestamp 1679581782
transform 1 0 11520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_121
timestamp 1679581782
transform 1 0 12192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_128
timestamp 1679581782
transform 1 0 12864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_135
timestamp 1679581782
transform 1 0 13536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_142
timestamp 1679581782
transform 1 0 14208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_149
timestamp 1679581782
transform 1 0 14880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_156
timestamp 1679581782
transform 1 0 15552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_163
timestamp 1679581782
transform 1 0 16224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_170
timestamp 1679581782
transform 1 0 16896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_177
timestamp 1679581782
transform 1 0 17568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_184
timestamp 1679581782
transform 1 0 18240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_191
timestamp 1679581782
transform 1 0 18912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_198
timestamp 1679581782
transform 1 0 19584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_205
timestamp 1679581782
transform 1 0 20256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_212
timestamp 1679581782
transform 1 0 20928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_219
timestamp 1679581782
transform 1 0 21600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_226
timestamp 1679581782
transform 1 0 22272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_233
timestamp 1679581782
transform 1 0 22944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_240
timestamp 1679581782
transform 1 0 23616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_247
timestamp 1679581782
transform 1 0 24288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_254
timestamp 1679581782
transform 1 0 24960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_261
timestamp 1679581782
transform 1 0 25632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_268
timestamp 1679581782
transform 1 0 26304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_275
timestamp 1679581782
transform 1 0 26976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_282
timestamp 1679581782
transform 1 0 27648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_289
timestamp 1679581782
transform 1 0 28320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_296
timestamp 1679581782
transform 1 0 28992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_303
timestamp 1679581782
transform 1 0 29664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_310
timestamp 1679581782
transform 1 0 30336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_317
timestamp 1679581782
transform 1 0 31008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_324
timestamp 1679581782
transform 1 0 31680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_331
timestamp 1679581782
transform 1 0 32352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_338
timestamp 1679581782
transform 1 0 33024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_345
timestamp 1679581782
transform 1 0 33696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_352
timestamp 1679581782
transform 1 0 34368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_359
timestamp 1679581782
transform 1 0 35040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_366
timestamp 1679581782
transform 1 0 35712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_373
timestamp 1679581782
transform 1 0 36384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_380
timestamp 1679581782
transform 1 0 37056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_387
timestamp 1679581782
transform 1 0 37728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_394
timestamp 1679581782
transform 1 0 38400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_401
timestamp 1679581782
transform 1 0 39072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_408
timestamp 1679581782
transform 1 0 39744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_415
timestamp 1679581782
transform 1 0 40416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_422
timestamp 1679581782
transform 1 0 41088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_429
timestamp 1679581782
transform 1 0 41760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_436
timestamp 1679581782
transform 1 0 42432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_443
timestamp 1679581782
transform 1 0 43104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_450
timestamp 1679581782
transform 1 0 43776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_457
timestamp 1679581782
transform 1 0 44448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_464
timestamp 1679581782
transform 1 0 45120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_471
timestamp 1679581782
transform 1 0 45792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_478
timestamp 1679581782
transform 1 0 46464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_485
timestamp 1679581782
transform 1 0 47136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_492
timestamp 1679581782
transform 1 0 47808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_499
timestamp 1679581782
transform 1 0 48480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_506
timestamp 1679581782
transform 1 0 49152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_513
timestamp 1679581782
transform 1 0 49824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_520
timestamp 1679581782
transform 1 0 50496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_527
timestamp 1679581782
transform 1 0 51168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_534
timestamp 1679581782
transform 1 0 51840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_541
timestamp 1679581782
transform 1 0 52512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_548
timestamp 1679581782
transform 1 0 53184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_559
timestamp 1679581782
transform 1 0 54240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_566
timestamp 1679581782
transform 1 0 54912 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_573
timestamp 1677579658
transform 1 0 55584 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_579
timestamp 1677579658
transform 1 0 56160 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_594
timestamp 1679581782
transform 1 0 57600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_601
timestamp 1679577901
transform 1 0 58272 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_605
timestamp 1677579658
transform 1 0 58656 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_639
timestamp 1677580104
transform 1 0 61920 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_645
timestamp 1679581782
transform 1 0 62496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_652
timestamp 1679577901
transform 1 0 63168 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_656
timestamp 1677579658
transform 1 0 63552 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_671
timestamp 1679581782
transform 1 0 64992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_678
timestamp 1679581782
transform 1 0 65664 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_685
timestamp 1677579658
transform 1 0 66336 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_697
timestamp 1679577901
transform 1 0 67488 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_701
timestamp 1677580104
transform 1 0 67872 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_775
timestamp 1679581782
transform 1 0 74976 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_782
timestamp 1677579658
transform 1 0 75648 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_810
timestamp 1679581782
transform 1 0 78336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_817
timestamp 1679577901
transform 1 0 79008 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_821
timestamp 1677580104
transform 1 0 79392 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_0
timestamp 1677580104
transform 1 0 576 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_2
timestamp 1677579658
transform 1 0 768 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_34
timestamp 1679577901
transform 1 0 3840 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 4608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 6624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 7968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 8640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 9984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 10656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 12672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 18720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679581782
transform 1 0 19392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679581782
transform 1 0 20064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679581782
transform 1 0 20736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679581782
transform 1 0 21408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679581782
transform 1 0 22080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679581782
transform 1 0 22752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679581782
transform 1 0 23424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679581782
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 27456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 28128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679581782
transform 1 0 28800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679581782
transform 1 0 29472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679581782
transform 1 0 30144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679581782
transform 1 0 30816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679581782
transform 1 0 31488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_329
timestamp 1679581782
transform 1 0 32160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_336
timestamp 1679581782
transform 1 0 32832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_343
timestamp 1679581782
transform 1 0 33504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679581782
transform 1 0 34176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679581782
transform 1 0 34848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679581782
transform 1 0 35520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679581782
transform 1 0 36192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679581782
transform 1 0 36864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679581782
transform 1 0 37536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679581782
transform 1 0 38208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679581782
transform 1 0 38880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679581782
transform 1 0 39552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679581782
transform 1 0 40224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679581782
transform 1 0 40896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679581782
transform 1 0 41568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679581782
transform 1 0 42240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679581782
transform 1 0 42912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_448
timestamp 1679581782
transform 1 0 43584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_455
timestamp 1679581782
transform 1 0 44256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_462
timestamp 1679581782
transform 1 0 44928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_469
timestamp 1679581782
transform 1 0 45600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_476
timestamp 1679581782
transform 1 0 46272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679581782
transform 1 0 46944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679581782
transform 1 0 47616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_497
timestamp 1679581782
transform 1 0 48288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_504
timestamp 1679581782
transform 1 0 48960 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_511
timestamp 1677580104
transform 1 0 49632 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_513
timestamp 1677579658
transform 1 0 49824 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_519
timestamp 1677579658
transform 1 0 50400 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_525
timestamp 1679577901
transform 1 0 50976 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_529
timestamp 1677579658
transform 1 0 51360 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_544
timestamp 1679581782
transform 1 0 52800 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_551
timestamp 1677580104
transform 1 0 53472 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_580
timestamp 1677580104
transform 1 0 56256 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_582
timestamp 1677579658
transform 1 0 56448 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_587
timestamp 1679581782
transform 1 0 56928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_594
timestamp 1679581782
transform 1 0 57600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_601
timestamp 1679581782
transform 1 0 58272 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_608
timestamp 1677580104
transform 1 0 58944 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_610
timestamp 1677579658
transform 1 0 59136 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_642
timestamp 1679581782
transform 1 0 62208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_649
timestamp 1679577901
transform 1 0 62880 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_657
timestamp 1677579658
transform 1 0 63648 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_668
timestamp 1679581782
transform 1 0 64704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_675
timestamp 1679581782
transform 1 0 65376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_687
timestamp 1679581782
transform 1 0 66528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_694
timestamp 1679581782
transform 1 0 67200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_701
timestamp 1679581782
transform 1 0 67872 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_718
timestamp 1677579658
transform 1 0 69504 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_724
timestamp 1679577901
transform 1 0 70080 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_728
timestamp 1677579658
transform 1 0 70464 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_756
timestamp 1679581782
transform 1 0 73152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_763
timestamp 1679581782
transform 1 0 73824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_770
timestamp 1679581782
transform 1 0 74496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_777
timestamp 1679577901
transform 1 0 75168 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_781
timestamp 1677580104
transform 1 0 75552 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_806
timestamp 1679581782
transform 1 0 77952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_813
timestamp 1679581782
transform 1 0 78624 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_820
timestamp 1677580104
transform 1 0 79296 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_822
timestamp 1677579658
transform 1 0 79488 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_8
timestamp 1679577901
transform 1 0 1344 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_16
timestamp 1677580104
transform 1 0 2112 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_28
timestamp 1677579658
transform 1 0 3264 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_75
timestamp 1679581782
transform 1 0 7776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_82
timestamp 1679581782
transform 1 0 8448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_89
timestamp 1679581782
transform 1 0 9120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_96
timestamp 1679581782
transform 1 0 9792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_103
timestamp 1679581782
transform 1 0 10464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_110
timestamp 1679581782
transform 1 0 11136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_117
timestamp 1679581782
transform 1 0 11808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_124
timestamp 1679581782
transform 1 0 12480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_131
timestamp 1679581782
transform 1 0 13152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_138
timestamp 1679581782
transform 1 0 13824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_145
timestamp 1679581782
transform 1 0 14496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_152
timestamp 1679581782
transform 1 0 15168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_159
timestamp 1679581782
transform 1 0 15840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_166
timestamp 1679581782
transform 1 0 16512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_173
timestamp 1679581782
transform 1 0 17184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_180
timestamp 1679581782
transform 1 0 17856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_187
timestamp 1679581782
transform 1 0 18528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_194
timestamp 1679581782
transform 1 0 19200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_201
timestamp 1679581782
transform 1 0 19872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_208
timestamp 1679581782
transform 1 0 20544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_215
timestamp 1679581782
transform 1 0 21216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_222
timestamp 1679581782
transform 1 0 21888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_229
timestamp 1679581782
transform 1 0 22560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_236
timestamp 1679581782
transform 1 0 23232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_243
timestamp 1679581782
transform 1 0 23904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_250
timestamp 1679581782
transform 1 0 24576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_257
timestamp 1679581782
transform 1 0 25248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_264
timestamp 1679581782
transform 1 0 25920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_271
timestamp 1679581782
transform 1 0 26592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_278
timestamp 1679581782
transform 1 0 27264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_285
timestamp 1679581782
transform 1 0 27936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_292
timestamp 1679581782
transform 1 0 28608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_299
timestamp 1679581782
transform 1 0 29280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_306
timestamp 1679581782
transform 1 0 29952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_313
timestamp 1679581782
transform 1 0 30624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_320
timestamp 1679581782
transform 1 0 31296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_327
timestamp 1679581782
transform 1 0 31968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_334
timestamp 1679581782
transform 1 0 32640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_341
timestamp 1679581782
transform 1 0 33312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_348
timestamp 1679581782
transform 1 0 33984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_355
timestamp 1679581782
transform 1 0 34656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_362
timestamp 1679581782
transform 1 0 35328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_369
timestamp 1679581782
transform 1 0 36000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_376
timestamp 1679581782
transform 1 0 36672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_383
timestamp 1679581782
transform 1 0 37344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_390
timestamp 1679581782
transform 1 0 38016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_397
timestamp 1679581782
transform 1 0 38688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_404
timestamp 1679581782
transform 1 0 39360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_411
timestamp 1679581782
transform 1 0 40032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_418
timestamp 1679581782
transform 1 0 40704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_425
timestamp 1679581782
transform 1 0 41376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_432
timestamp 1679581782
transform 1 0 42048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_439
timestamp 1679581782
transform 1 0 42720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_446
timestamp 1679581782
transform 1 0 43392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_453
timestamp 1679581782
transform 1 0 44064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_460
timestamp 1679581782
transform 1 0 44736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_467
timestamp 1679581782
transform 1 0 45408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_474
timestamp 1679581782
transform 1 0 46080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_481
timestamp 1679577901
transform 1 0 46752 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_485
timestamp 1677580104
transform 1 0 47136 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_492
timestamp 1679581782
transform 1 0 47808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_499
timestamp 1679581782
transform 1 0 48480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_506
timestamp 1679577901
transform 1 0 49152 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_537
timestamp 1677579658
transform 1 0 52128 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_569
timestamp 1677580104
transform 1 0 55200 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_571
timestamp 1677579658
transform 1 0 55392 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_592
timestamp 1679577901
transform 1 0 57408 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_596
timestamp 1677579658
transform 1 0 57792 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_602
timestamp 1679577901
transform 1 0 58368 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_606
timestamp 1677579658
transform 1 0 58752 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_612
timestamp 1679581782
transform 1 0 59328 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_619
timestamp 1677579658
transform 1 0 60000 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_624
timestamp 1679581782
transform 1 0 60480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_631
timestamp 1679581782
transform 1 0 61152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_638
timestamp 1679581782
transform 1 0 61824 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_645
timestamp 1677580104
transform 1 0 62496 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_647
timestamp 1677579658
transform 1 0 62688 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_739
timestamp 1677580104
transform 1 0 71520 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_741
timestamp 1677579658
transform 1 0 71712 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_4
timestamp 1677580104
transform 1 0 960 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_20
timestamp 1679581782
transform 1 0 2496 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_27
timestamp 1677580104
transform 1 0 3168 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_50
timestamp 1677579658
transform 1 0 5376 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_59
timestamp 1679581782
transform 1 0 6240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_66
timestamp 1679581782
transform 1 0 6912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_73
timestamp 1679581782
transform 1 0 7584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_80
timestamp 1679581782
transform 1 0 8256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_87
timestamp 1679581782
transform 1 0 8928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_94
timestamp 1679581782
transform 1 0 9600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_101
timestamp 1679581782
transform 1 0 10272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_108
timestamp 1679581782
transform 1 0 10944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_115
timestamp 1679581782
transform 1 0 11616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_122
timestamp 1679581782
transform 1 0 12288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_129
timestamp 1679581782
transform 1 0 12960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_136
timestamp 1679581782
transform 1 0 13632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_143
timestamp 1679581782
transform 1 0 14304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_150
timestamp 1679581782
transform 1 0 14976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_157
timestamp 1679581782
transform 1 0 15648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_164
timestamp 1679581782
transform 1 0 16320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_171
timestamp 1679581782
transform 1 0 16992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_178
timestamp 1679581782
transform 1 0 17664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_185
timestamp 1679581782
transform 1 0 18336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_192
timestamp 1679581782
transform 1 0 19008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_199
timestamp 1679581782
transform 1 0 19680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_206
timestamp 1679581782
transform 1 0 20352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_213
timestamp 1679581782
transform 1 0 21024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_220
timestamp 1679581782
transform 1 0 21696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_227
timestamp 1679581782
transform 1 0 22368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_234
timestamp 1679581782
transform 1 0 23040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_241
timestamp 1679581782
transform 1 0 23712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_248
timestamp 1679581782
transform 1 0 24384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_255
timestamp 1679581782
transform 1 0 25056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_262
timestamp 1679581782
transform 1 0 25728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_269
timestamp 1679581782
transform 1 0 26400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_276
timestamp 1679581782
transform 1 0 27072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_283
timestamp 1679581782
transform 1 0 27744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_290
timestamp 1679581782
transform 1 0 28416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_297
timestamp 1679581782
transform 1 0 29088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_304
timestamp 1679581782
transform 1 0 29760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_311
timestamp 1679581782
transform 1 0 30432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_318
timestamp 1679581782
transform 1 0 31104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_325
timestamp 1679581782
transform 1 0 31776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_332
timestamp 1679581782
transform 1 0 32448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_339
timestamp 1679581782
transform 1 0 33120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_346
timestamp 1679581782
transform 1 0 33792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_353
timestamp 1679581782
transform 1 0 34464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_360
timestamp 1679581782
transform 1 0 35136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_367
timestamp 1679581782
transform 1 0 35808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_374
timestamp 1679581782
transform 1 0 36480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_381
timestamp 1679581782
transform 1 0 37152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_388
timestamp 1679581782
transform 1 0 37824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_395
timestamp 1679581782
transform 1 0 38496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_402
timestamp 1679581782
transform 1 0 39168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_409
timestamp 1679581782
transform 1 0 39840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_416
timestamp 1679581782
transform 1 0 40512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_423
timestamp 1679581782
transform 1 0 41184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_430
timestamp 1679581782
transform 1 0 41856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_437
timestamp 1679581782
transform 1 0 42528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_444
timestamp 1679581782
transform 1 0 43200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_451
timestamp 1679581782
transform 1 0 43872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_458
timestamp 1679581782
transform 1 0 44544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_465
timestamp 1679577901
transform 1 0 45216 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_496
timestamp 1677580104
transform 1 0 48192 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_507
timestamp 1679581782
transform 1 0 49248 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_514
timestamp 1677579658
transform 1 0 49920 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_519
timestamp 1679581782
transform 1 0 50400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_526
timestamp 1679577901
transform 1 0 51072 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_548
timestamp 1679581782
transform 1 0 53184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_555
timestamp 1679581782
transform 1 0 53856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_562
timestamp 1679581782
transform 1 0 54528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_569
timestamp 1679577901
transform 1 0 55200 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_605
timestamp 1677579658
transform 1 0 58656 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_648
timestamp 1677579658
transform 1 0 62784 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_681
timestamp 1677579658
transform 1 0 65952 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_694
timestamp 1679581782
transform 1 0 67200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_701
timestamp 1679581782
transform 1 0 67872 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_708
timestamp 1677580104
transform 1 0 68544 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_719
timestamp 1679581782
transform 1 0 69600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_726
timestamp 1679581782
transform 1 0 70272 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_733
timestamp 1677580104
transform 1 0 70944 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_744
timestamp 1677580104
transform 1 0 72000 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_746
timestamp 1677579658
transform 1 0 72192 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_751
timestamp 1679581782
transform 1 0 72672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_758
timestamp 1679581782
transform 1 0 73344 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_765
timestamp 1677580104
transform 1 0 74016 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_771
timestamp 1679581782
transform 1 0 74592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_778
timestamp 1679577901
transform 1 0 75264 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_782
timestamp 1677580104
transform 1 0 75648 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_794
timestamp 1677580104
transform 1 0 76800 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_796
timestamp 1677579658
transform 1 0 76992 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_802
timestamp 1677580104
transform 1 0 77568 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679581782
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679581782
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_822
timestamp 1677579658
transform 1 0 79488 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 576 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_33
timestamp 1679577901
transform 1 0 3744 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_61
timestamp 1679581782
transform 1 0 6432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_68
timestamp 1679581782
transform 1 0 7104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_75
timestamp 1679581782
transform 1 0 7776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_82
timestamp 1679581782
transform 1 0 8448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_89
timestamp 1679581782
transform 1 0 9120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_96
timestamp 1679581782
transform 1 0 9792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_103
timestamp 1679581782
transform 1 0 10464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_110
timestamp 1679581782
transform 1 0 11136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_117
timestamp 1679581782
transform 1 0 11808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_124
timestamp 1679581782
transform 1 0 12480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_131
timestamp 1679581782
transform 1 0 13152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_138
timestamp 1679581782
transform 1 0 13824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_145
timestamp 1679581782
transform 1 0 14496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_152
timestamp 1679581782
transform 1 0 15168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_159
timestamp 1679581782
transform 1 0 15840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_166
timestamp 1679581782
transform 1 0 16512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_173
timestamp 1679581782
transform 1 0 17184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_180
timestamp 1679581782
transform 1 0 17856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_187
timestamp 1679581782
transform 1 0 18528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_194
timestamp 1679581782
transform 1 0 19200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_201
timestamp 1679581782
transform 1 0 19872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_208
timestamp 1679581782
transform 1 0 20544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_215
timestamp 1679581782
transform 1 0 21216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_222
timestamp 1679581782
transform 1 0 21888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_229
timestamp 1679581782
transform 1 0 22560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_236
timestamp 1679581782
transform 1 0 23232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_243
timestamp 1679581782
transform 1 0 23904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_250
timestamp 1679581782
transform 1 0 24576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_257
timestamp 1679581782
transform 1 0 25248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_264
timestamp 1679581782
transform 1 0 25920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_271
timestamp 1679581782
transform 1 0 26592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_278
timestamp 1679581782
transform 1 0 27264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_285
timestamp 1679581782
transform 1 0 27936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_292
timestamp 1679581782
transform 1 0 28608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_299
timestamp 1679581782
transform 1 0 29280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_306
timestamp 1679581782
transform 1 0 29952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_313
timestamp 1679581782
transform 1 0 30624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_320
timestamp 1679581782
transform 1 0 31296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_327
timestamp 1679581782
transform 1 0 31968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_334
timestamp 1679581782
transform 1 0 32640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_341
timestamp 1679581782
transform 1 0 33312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_348
timestamp 1679581782
transform 1 0 33984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_355
timestamp 1679581782
transform 1 0 34656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_362
timestamp 1679581782
transform 1 0 35328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_369
timestamp 1679581782
transform 1 0 36000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_376
timestamp 1679581782
transform 1 0 36672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_383
timestamp 1679581782
transform 1 0 37344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_390
timestamp 1679581782
transform 1 0 38016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_397
timestamp 1679581782
transform 1 0 38688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_404
timestamp 1679581782
transform 1 0 39360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_411
timestamp 1679581782
transform 1 0 40032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_418
timestamp 1679581782
transform 1 0 40704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_425
timestamp 1679581782
transform 1 0 41376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_432
timestamp 1679581782
transform 1 0 42048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_439
timestamp 1679581782
transform 1 0 42720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_446
timestamp 1679581782
transform 1 0 43392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_453
timestamp 1679581782
transform 1 0 44064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_460
timestamp 1679581782
transform 1 0 44736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_467
timestamp 1679581782
transform 1 0 45408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_478
timestamp 1679581782
transform 1 0 46464 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_490
timestamp 1677580104
transform 1 0 47616 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_492
timestamp 1677579658
transform 1 0 47808 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_512
timestamp 1679581782
transform 1 0 49728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_519
timestamp 1679581782
transform 1 0 50400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_526
timestamp 1679581782
transform 1 0 51072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_533
timestamp 1679577901
transform 1 0 51744 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_547
timestamp 1679577901
transform 1 0 53088 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_551
timestamp 1677580104
transform 1 0 53472 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_567
timestamp 1679581782
transform 1 0 55008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_574
timestamp 1679577901
transform 1 0 55680 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_578
timestamp 1677579658
transform 1 0 56064 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_587
timestamp 1679581782
transform 1 0 56928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_594
timestamp 1679581782
transform 1 0 57600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_601
timestamp 1679581782
transform 1 0 58272 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_608
timestamp 1677580104
transform 1 0 58944 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_619
timestamp 1677580104
transform 1 0 60000 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_658
timestamp 1679581782
transform 1 0 63744 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_665
timestamp 1677579658
transform 1 0 64416 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679581782
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_683
timestamp 1677579658
transform 1 0 66144 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_689
timestamp 1679577901
transform 1 0 66720 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679581782
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679581782
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_711
timestamp 1679577901
transform 1 0 68832 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679581782
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_732
timestamp 1677580104
transform 1 0 70848 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_734
timestamp 1677579658
transform 1 0 71040 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_753
timestamp 1679581782
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_792
timestamp 1679577901
transform 1 0 76608 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_796
timestamp 1677579658
transform 1 0 76992 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_802
timestamp 1679581782
transform 1 0 77568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_809
timestamp 1679581782
transform 1 0 78240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679581782
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_7
timestamp 1679577901
transform 1 0 1248 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679581782
transform 1 0 2976 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_32
timestamp 1677579658
transform 1 0 3648 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_43
timestamp 1677580104
transform 1 0 4704 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_45
timestamp 1677579658
transform 1 0 4896 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_73
timestamp 1679581782
transform 1 0 7584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_80
timestamp 1679581782
transform 1 0 8256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_87
timestamp 1679581782
transform 1 0 8928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_94
timestamp 1679581782
transform 1 0 9600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_101
timestamp 1679581782
transform 1 0 10272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_108
timestamp 1679581782
transform 1 0 10944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_115
timestamp 1679581782
transform 1 0 11616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_122
timestamp 1679581782
transform 1 0 12288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_129
timestamp 1679581782
transform 1 0 12960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_136
timestamp 1679581782
transform 1 0 13632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_143
timestamp 1679581782
transform 1 0 14304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_150
timestamp 1679581782
transform 1 0 14976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_157
timestamp 1679581782
transform 1 0 15648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_164
timestamp 1679581782
transform 1 0 16320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_171
timestamp 1679581782
transform 1 0 16992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_178
timestamp 1679581782
transform 1 0 17664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_185
timestamp 1679581782
transform 1 0 18336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_192
timestamp 1679581782
transform 1 0 19008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_199
timestamp 1679581782
transform 1 0 19680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_206
timestamp 1679581782
transform 1 0 20352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_213
timestamp 1679581782
transform 1 0 21024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_220
timestamp 1679581782
transform 1 0 21696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_227
timestamp 1679581782
transform 1 0 22368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_234
timestamp 1679581782
transform 1 0 23040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_241
timestamp 1679581782
transform 1 0 23712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_248
timestamp 1679581782
transform 1 0 24384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_255
timestamp 1679581782
transform 1 0 25056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_262
timestamp 1679581782
transform 1 0 25728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_269
timestamp 1679581782
transform 1 0 26400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_276
timestamp 1679581782
transform 1 0 27072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_283
timestamp 1679581782
transform 1 0 27744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_290
timestamp 1679581782
transform 1 0 28416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_297
timestamp 1679581782
transform 1 0 29088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_304
timestamp 1679581782
transform 1 0 29760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_311
timestamp 1679581782
transform 1 0 30432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_318
timestamp 1679581782
transform 1 0 31104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_325
timestamp 1679581782
transform 1 0 31776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_332
timestamp 1679581782
transform 1 0 32448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_339
timestamp 1679581782
transform 1 0 33120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_346
timestamp 1679581782
transform 1 0 33792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_353
timestamp 1679581782
transform 1 0 34464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_360
timestamp 1679581782
transform 1 0 35136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_367
timestamp 1679581782
transform 1 0 35808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_374
timestamp 1679581782
transform 1 0 36480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_381
timestamp 1679581782
transform 1 0 37152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_388
timestamp 1679581782
transform 1 0 37824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_395
timestamp 1679581782
transform 1 0 38496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_402
timestamp 1679581782
transform 1 0 39168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_409
timestamp 1679581782
transform 1 0 39840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_416
timestamp 1679581782
transform 1 0 40512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_423
timestamp 1679581782
transform 1 0 41184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_430
timestamp 1679581782
transform 1 0 41856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_437
timestamp 1679581782
transform 1 0 42528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_444
timestamp 1679581782
transform 1 0 43200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_451
timestamp 1679581782
transform 1 0 43872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_458
timestamp 1679581782
transform 1 0 44544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_465
timestamp 1679581782
transform 1 0 45216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_472
timestamp 1679581782
transform 1 0 45888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_479
timestamp 1679577901
transform 1 0 46560 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_483
timestamp 1677580104
transform 1 0 46944 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_495
timestamp 1677580104
transform 1 0 48096 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_501
timestamp 1677579658
transform 1 0 48672 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_556
timestamp 1677579658
transform 1 0 53952 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_589
timestamp 1677579658
transform 1 0 57120 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_594
timestamp 1679577901
transform 1 0 57600 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_608
timestamp 1677580104
transform 1 0 58944 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_615
timestamp 1679577901
transform 1 0 59616 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_619
timestamp 1677579658
transform 1 0 60000 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_624
timestamp 1679577901
transform 1 0 60480 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_628
timestamp 1677579658
transform 1 0 60864 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_634
timestamp 1677580104
transform 1 0 61440 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_640
timestamp 1679581782
transform 1 0 62016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_647
timestamp 1679581782
transform 1 0 62688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_658
timestamp 1679581782
transform 1 0 63744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_665
timestamp 1679581782
transform 1 0 64416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_672
timestamp 1679577901
transform 1 0 65088 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_686
timestamp 1677579658
transform 1 0 66432 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_741
timestamp 1677580104
transform 1 0 71712 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_774
timestamp 1679581782
transform 1 0 74880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_4
timestamp 1679577901
transform 1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_8
timestamp 1677579658
transform 1 0 1344 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_36
timestamp 1677579658
transform 1 0 4032 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_41
timestamp 1679577901
transform 1 0 4512 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_49
timestamp 1677580104
transform 1 0 5280 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_55
timestamp 1679581782
transform 1 0 5856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_62
timestamp 1679581782
transform 1 0 6528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_69
timestamp 1679581782
transform 1 0 7200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_76
timestamp 1679581782
transform 1 0 7872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_83
timestamp 1679581782
transform 1 0 8544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_90
timestamp 1679581782
transform 1 0 9216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_97
timestamp 1679581782
transform 1 0 9888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_104
timestamp 1679581782
transform 1 0 10560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_111
timestamp 1679581782
transform 1 0 11232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_118
timestamp 1679581782
transform 1 0 11904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_125
timestamp 1679581782
transform 1 0 12576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_132
timestamp 1679581782
transform 1 0 13248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_139
timestamp 1679581782
transform 1 0 13920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_146
timestamp 1679581782
transform 1 0 14592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_153
timestamp 1679581782
transform 1 0 15264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_160
timestamp 1679581782
transform 1 0 15936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_167
timestamp 1679581782
transform 1 0 16608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_174
timestamp 1679581782
transform 1 0 17280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_181
timestamp 1679581782
transform 1 0 17952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_188
timestamp 1679581782
transform 1 0 18624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_195
timestamp 1679581782
transform 1 0 19296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_202
timestamp 1679581782
transform 1 0 19968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_209
timestamp 1679581782
transform 1 0 20640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_216
timestamp 1679581782
transform 1 0 21312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_223
timestamp 1679581782
transform 1 0 21984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_230
timestamp 1679581782
transform 1 0 22656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_237
timestamp 1679581782
transform 1 0 23328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_244
timestamp 1679581782
transform 1 0 24000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_251
timestamp 1679581782
transform 1 0 24672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_258
timestamp 1679581782
transform 1 0 25344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_265
timestamp 1679581782
transform 1 0 26016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_272
timestamp 1679581782
transform 1 0 26688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_279
timestamp 1679581782
transform 1 0 27360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_286
timestamp 1679581782
transform 1 0 28032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_293
timestamp 1679581782
transform 1 0 28704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_300
timestamp 1679581782
transform 1 0 29376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_307
timestamp 1679581782
transform 1 0 30048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_314
timestamp 1679581782
transform 1 0 30720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_321
timestamp 1679581782
transform 1 0 31392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_328
timestamp 1679581782
transform 1 0 32064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_335
timestamp 1679581782
transform 1 0 32736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_342
timestamp 1679581782
transform 1 0 33408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_349
timestamp 1679581782
transform 1 0 34080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_356
timestamp 1679581782
transform 1 0 34752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_363
timestamp 1679581782
transform 1 0 35424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_370
timestamp 1679581782
transform 1 0 36096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_377
timestamp 1679581782
transform 1 0 36768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_384
timestamp 1679581782
transform 1 0 37440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_391
timestamp 1679581782
transform 1 0 38112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_398
timestamp 1679581782
transform 1 0 38784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_405
timestamp 1679581782
transform 1 0 39456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_412
timestamp 1679581782
transform 1 0 40128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_419
timestamp 1679581782
transform 1 0 40800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_426
timestamp 1679581782
transform 1 0 41472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_433
timestamp 1679581782
transform 1 0 42144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_440
timestamp 1679581782
transform 1 0 42816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_447
timestamp 1679581782
transform 1 0 43488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_454
timestamp 1679581782
transform 1 0 44160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_461
timestamp 1679577901
transform 1 0 44832 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_465
timestamp 1677579658
transform 1 0 45216 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_493
timestamp 1679581782
transform 1 0 47904 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_500
timestamp 1677579658
transform 1 0 48576 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_528
timestamp 1679577901
transform 1 0 51264 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_532
timestamp 1677580104
transform 1 0 51648 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_538
timestamp 1679577901
transform 1 0 52224 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_542
timestamp 1677579658
transform 1 0 52608 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_553
timestamp 1679577901
transform 1 0 53664 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_557
timestamp 1677580104
transform 1 0 54048 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_571
timestamp 1679581782
transform 1 0 55392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_578
timestamp 1679581782
transform 1 0 56064 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_612
timestamp 1677580104
transform 1 0 59328 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_629
timestamp 1679581782
transform 1 0 60960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_636
timestamp 1679577901
transform 1 0 61632 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_640
timestamp 1677579658
transform 1 0 62016 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_677
timestamp 1677580104
transform 1 0 65568 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_691
timestamp 1679581782
transform 1 0 66912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_698
timestamp 1679581782
transform 1 0 67584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_705
timestamp 1679581782
transform 1 0 68256 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_712
timestamp 1677580104
transform 1 0 68928 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 70464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_735
timestamp 1679577901
transform 1 0 71136 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_739
timestamp 1677579658
transform 1 0 71520 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_745
timestamp 1677580104
transform 1 0 72096 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_747
timestamp 1677579658
transform 1 0 72288 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_752
timestamp 1679581782
transform 1 0 72768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_759
timestamp 1679581782
transform 1 0 73440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_766
timestamp 1679581782
transform 1 0 74112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_773
timestamp 1679581782
transform 1 0 74784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_790
timestamp 1679577901
transform 1 0 76416 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_794
timestamp 1677579658
transform 1 0 76800 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_799
timestamp 1677579658
transform 1 0 77280 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_808
timestamp 1679581782
transform 1 0 78144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_815
timestamp 1679581782
transform 1 0 78816 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_822
timestamp 1677579658
transform 1 0 79488 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_27
timestamp 1677579658
transform 1 0 3168 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_38
timestamp 1677580104
transform 1 0 4224 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_40
timestamp 1677579658
transform 1 0 4416 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_73
timestamp 1679581782
transform 1 0 7584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_80
timestamp 1679581782
transform 1 0 8256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_87
timestamp 1679581782
transform 1 0 8928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_94
timestamp 1679581782
transform 1 0 9600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_101
timestamp 1679581782
transform 1 0 10272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_108
timestamp 1679581782
transform 1 0 10944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_115
timestamp 1679581782
transform 1 0 11616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_122
timestamp 1679581782
transform 1 0 12288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_129
timestamp 1679581782
transform 1 0 12960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_136
timestamp 1679581782
transform 1 0 13632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_143
timestamp 1679581782
transform 1 0 14304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_150
timestamp 1679581782
transform 1 0 14976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_157
timestamp 1679581782
transform 1 0 15648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_164
timestamp 1679581782
transform 1 0 16320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_171
timestamp 1679581782
transform 1 0 16992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_178
timestamp 1679581782
transform 1 0 17664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_185
timestamp 1679581782
transform 1 0 18336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_192
timestamp 1679581782
transform 1 0 19008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_199
timestamp 1679581782
transform 1 0 19680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_206
timestamp 1679581782
transform 1 0 20352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_213
timestamp 1679581782
transform 1 0 21024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_220
timestamp 1679581782
transform 1 0 21696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_227
timestamp 1679581782
transform 1 0 22368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_234
timestamp 1679581782
transform 1 0 23040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_241
timestamp 1679581782
transform 1 0 23712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_248
timestamp 1679581782
transform 1 0 24384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_255
timestamp 1679581782
transform 1 0 25056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_262
timestamp 1679581782
transform 1 0 25728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_269
timestamp 1679581782
transform 1 0 26400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_276
timestamp 1679581782
transform 1 0 27072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_283
timestamp 1679581782
transform 1 0 27744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_290
timestamp 1679581782
transform 1 0 28416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_297
timestamp 1679581782
transform 1 0 29088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_304
timestamp 1679581782
transform 1 0 29760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_311
timestamp 1679581782
transform 1 0 30432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_318
timestamp 1679581782
transform 1 0 31104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_325
timestamp 1679581782
transform 1 0 31776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_332
timestamp 1679581782
transform 1 0 32448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_339
timestamp 1679581782
transform 1 0 33120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_346
timestamp 1679581782
transform 1 0 33792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_353
timestamp 1679581782
transform 1 0 34464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_360
timestamp 1679581782
transform 1 0 35136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_367
timestamp 1679581782
transform 1 0 35808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_374
timestamp 1679581782
transform 1 0 36480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_381
timestamp 1679581782
transform 1 0 37152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_388
timestamp 1679581782
transform 1 0 37824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_395
timestamp 1679581782
transform 1 0 38496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_402
timestamp 1679581782
transform 1 0 39168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_409
timestamp 1679581782
transform 1 0 39840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_416
timestamp 1679581782
transform 1 0 40512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_423
timestamp 1679581782
transform 1 0 41184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_430
timestamp 1679581782
transform 1 0 41856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_437
timestamp 1679581782
transform 1 0 42528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_444
timestamp 1679581782
transform 1 0 43200 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_451
timestamp 1677580104
transform 1 0 43872 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_458
timestamp 1677580104
transform 1 0 44544 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_465
timestamp 1677579658
transform 1 0 45216 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_475
timestamp 1679577901
transform 1 0 46176 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_479
timestamp 1677579658
transform 1 0 46560 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_490
timestamp 1677580104
transform 1 0 47616 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_551
timestamp 1679577901
transform 1 0 53472 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_555
timestamp 1677579658
transform 1 0 53856 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_561
timestamp 1679581782
transform 1 0 54432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_568
timestamp 1679581782
transform 1 0 55104 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_575
timestamp 1677579658
transform 1 0 55776 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_608
timestamp 1679581782
transform 1 0 58944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_615
timestamp 1679577901
transform 1 0 59616 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_654
timestamp 1677580104
transform 1 0 63360 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_735
timestamp 1677580104
transform 1 0 71136 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679581782
transform 1 0 71808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679581782
transform 1 0 72480 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_756
timestamp 1677580104
transform 1 0 73152 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_758
timestamp 1677579658
transform 1 0 73344 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_800
timestamp 1677580104
transform 1 0 77376 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_802
timestamp 1677579658
transform 1 0 77568 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679581782
transform 1 0 78048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679581782
transform 1 0 78720 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_821
timestamp 1677580104
transform 1 0 79392 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_4
timestamp 1677579658
transform 1 0 960 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_39
timestamp 1679577901
transform 1 0 4320 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_47
timestamp 1679581782
transform 1 0 5088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_54
timestamp 1679581782
transform 1 0 5760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_61
timestamp 1679581782
transform 1 0 6432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_68
timestamp 1679581782
transform 1 0 7104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_75
timestamp 1679581782
transform 1 0 7776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_82
timestamp 1679581782
transform 1 0 8448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_89
timestamp 1679581782
transform 1 0 9120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_96
timestamp 1679581782
transform 1 0 9792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_103
timestamp 1679581782
transform 1 0 10464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_110
timestamp 1679581782
transform 1 0 11136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_117
timestamp 1679581782
transform 1 0 11808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_124
timestamp 1679581782
transform 1 0 12480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_131
timestamp 1679581782
transform 1 0 13152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_138
timestamp 1679581782
transform 1 0 13824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_145
timestamp 1679581782
transform 1 0 14496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_152
timestamp 1679581782
transform 1 0 15168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_159
timestamp 1679581782
transform 1 0 15840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_166
timestamp 1679581782
transform 1 0 16512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_173
timestamp 1679581782
transform 1 0 17184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_180
timestamp 1679581782
transform 1 0 17856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_187
timestamp 1679581782
transform 1 0 18528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_194
timestamp 1679581782
transform 1 0 19200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_201
timestamp 1679581782
transform 1 0 19872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_208
timestamp 1679581782
transform 1 0 20544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_215
timestamp 1679581782
transform 1 0 21216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_222
timestamp 1679581782
transform 1 0 21888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_229
timestamp 1679581782
transform 1 0 22560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_236
timestamp 1679581782
transform 1 0 23232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_243
timestamp 1679581782
transform 1 0 23904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_250
timestamp 1679581782
transform 1 0 24576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_257
timestamp 1679581782
transform 1 0 25248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_264
timestamp 1679581782
transform 1 0 25920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_271
timestamp 1679581782
transform 1 0 26592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_278
timestamp 1679581782
transform 1 0 27264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_285
timestamp 1679581782
transform 1 0 27936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_292
timestamp 1679581782
transform 1 0 28608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_299
timestamp 1679581782
transform 1 0 29280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_306
timestamp 1679581782
transform 1 0 29952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_313
timestamp 1679581782
transform 1 0 30624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_320
timestamp 1679581782
transform 1 0 31296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_327
timestamp 1679581782
transform 1 0 31968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_334
timestamp 1679581782
transform 1 0 32640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_341
timestamp 1679581782
transform 1 0 33312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_348
timestamp 1679581782
transform 1 0 33984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_355
timestamp 1679581782
transform 1 0 34656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_362
timestamp 1679581782
transform 1 0 35328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_369
timestamp 1679581782
transform 1 0 36000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_376
timestamp 1679581782
transform 1 0 36672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_383
timestamp 1679581782
transform 1 0 37344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_390
timestamp 1679581782
transform 1 0 38016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_397
timestamp 1679581782
transform 1 0 38688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_404
timestamp 1679581782
transform 1 0 39360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_411
timestamp 1679581782
transform 1 0 40032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_418
timestamp 1679581782
transform 1 0 40704 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_425
timestamp 1677579658
transform 1 0 41376 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_453
timestamp 1677579658
transform 1 0 44064 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_481
timestamp 1679581782
transform 1 0 46752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_488
timestamp 1679581782
transform 1 0 47424 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_495
timestamp 1677580104
transform 1 0 48096 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_497
timestamp 1677579658
transform 1 0 48288 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679581782
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_522
timestamp 1677580104
transform 1 0 50688 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_533
timestamp 1679577901
transform 1 0 51744 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_557
timestamp 1677580104
transform 1 0 54048 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_559
timestamp 1677579658
transform 1 0 54240 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_587
timestamp 1679581782
transform 1 0 56928 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_594
timestamp 1677579658
transform 1 0 57600 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_604
timestamp 1677579658
transform 1 0 58560 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_622
timestamp 1679577901
transform 1 0 60288 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_626
timestamp 1677580104
transform 1 0 60672 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_632
timestamp 1679581782
transform 1 0 61248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_639
timestamp 1679581782
transform 1 0 61920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_646
timestamp 1679581782
transform 1 0 62592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_653
timestamp 1679577901
transform 1 0 63264 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_657
timestamp 1677579658
transform 1 0 63648 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_672
timestamp 1679581782
transform 1 0 65088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_679
timestamp 1679581782
transform 1 0 65760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679581782
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679581782
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_704
timestamp 1677579658
transform 1 0 68160 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_727
timestamp 1677580104
transform 1 0 70368 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_729
timestamp 1677579658
transform 1 0 70560 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_771
timestamp 1679581782
transform 1 0 74592 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_778
timestamp 1677580104
transform 1 0 75264 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_780
timestamp 1677579658
transform 1 0 75456 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_4
timestamp 1677579658
transform 1 0 960 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_13
timestamp 1677579658
transform 1 0 1824 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_19
timestamp 1677580104
transform 1 0 2400 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_21
timestamp 1677579658
transform 1 0 2592 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_36
timestamp 1677580104
transform 1 0 4032 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679581782
transform 1 0 7296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679581782
transform 1 0 7968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679581782
transform 1 0 8640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679581782
transform 1 0 9312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679581782
transform 1 0 9984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 10656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 11328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679581782
transform 1 0 12000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679581782
transform 1 0 12672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679581782
transform 1 0 13344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679581782
transform 1 0 14016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679581782
transform 1 0 14688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679581782
transform 1 0 15360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679581782
transform 1 0 16032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679581782
transform 1 0 16704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679581782
transform 1 0 17376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679581782
transform 1 0 18048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 18720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679581782
transform 1 0 19392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_203
timestamp 1679581782
transform 1 0 20064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_210
timestamp 1679581782
transform 1 0 20736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679581782
transform 1 0 21408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679581782
transform 1 0 22080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679581782
transform 1 0 22752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679581782
transform 1 0 23424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_245
timestamp 1679581782
transform 1 0 24096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_252
timestamp 1679581782
transform 1 0 24768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_259
timestamp 1679581782
transform 1 0 25440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_266
timestamp 1679581782
transform 1 0 26112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679581782
transform 1 0 26784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679581782
transform 1 0 27456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1679581782
transform 1 0 28128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1679581782
transform 1 0 28800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1679581782
transform 1 0 29472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1679581782
transform 1 0 30144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679581782
transform 1 0 30816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_322
timestamp 1679581782
transform 1 0 31488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_329
timestamp 1679581782
transform 1 0 32160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_336
timestamp 1679581782
transform 1 0 32832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679581782
transform 1 0 33504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679581782
transform 1 0 34176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_357
timestamp 1679581782
transform 1 0 34848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_364
timestamp 1679581782
transform 1 0 35520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_371
timestamp 1679581782
transform 1 0 36192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_378
timestamp 1679581782
transform 1 0 36864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_385
timestamp 1679581782
transform 1 0 37536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_392
timestamp 1679581782
transform 1 0 38208 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_399
timestamp 1677580104
transform 1 0 38880 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_406
timestamp 1677580104
transform 1 0 39552 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_408
timestamp 1677579658
transform 1 0 39744 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_414
timestamp 1677580104
transform 1 0 40320 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_421
timestamp 1677580104
transform 1 0 40992 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_442
timestamp 1679581782
transform 1 0 43008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_449
timestamp 1679581782
transform 1 0 43680 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_456
timestamp 1677580104
transform 1 0 44352 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_458
timestamp 1677579658
transform 1 0 44544 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_463
timestamp 1679581782
transform 1 0 45024 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_470
timestamp 1677579658
transform 1 0 45696 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_489
timestamp 1679581782
transform 1 0 47520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_496
timestamp 1679581782
transform 1 0 48192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_503
timestamp 1679581782
transform 1 0 48864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_510
timestamp 1679577901
transform 1 0 49536 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_514
timestamp 1677580104
transform 1 0 49920 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_550
timestamp 1677580104
transform 1 0 53376 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_552
timestamp 1677579658
transform 1 0 53568 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_557
timestamp 1677579658
transform 1 0 54048 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_562
timestamp 1677580104
transform 1 0 54528 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_564
timestamp 1677579658
transform 1 0 54720 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_569
timestamp 1679581782
transform 1 0 55200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_576
timestamp 1679577901
transform 1 0 55872 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_580
timestamp 1677579658
transform 1 0 56256 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_585
timestamp 1679577901
transform 1 0 56736 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_589
timestamp 1677580104
transform 1 0 57120 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_677
timestamp 1679581782
transform 1 0 65568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_684
timestamp 1679577901
transform 1 0 66240 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_688
timestamp 1677580104
transform 1 0 66624 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_734
timestamp 1677580104
transform 1 0 71040 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_744
timestamp 1677579658
transform 1 0 72000 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679581782
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679581782
transform 1 0 73152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_767
timestamp 1679581782
transform 1 0 74208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_774
timestamp 1679577901
transform 1 0 74880 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_778
timestamp 1677580104
transform 1 0 75264 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_794
timestamp 1677580104
transform 1 0 76800 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_809
timestamp 1679581782
transform 1 0 78240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_816
timestamp 1679581782
transform 1 0 78912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_4
timestamp 1679577901
transform 1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_8
timestamp 1677579658
transform 1 0 1344 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_13
timestamp 1677580104
transform 1 0 1824 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_15
timestamp 1677579658
transform 1 0 2016 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_30
timestamp 1679581782
transform 1 0 3456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_37
timestamp 1679581782
transform 1 0 4128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_44
timestamp 1679577901
transform 1 0 4800 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_52
timestamp 1679581782
transform 1 0 5568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_59
timestamp 1679581782
transform 1 0 6240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_66
timestamp 1679581782
transform 1 0 6912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_73
timestamp 1679581782
transform 1 0 7584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_80
timestamp 1679581782
transform 1 0 8256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_87
timestamp 1679581782
transform 1 0 8928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_94
timestamp 1679581782
transform 1 0 9600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_101
timestamp 1679581782
transform 1 0 10272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_108
timestamp 1679581782
transform 1 0 10944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_115
timestamp 1679581782
transform 1 0 11616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_122
timestamp 1679581782
transform 1 0 12288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_129
timestamp 1679581782
transform 1 0 12960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_136
timestamp 1679581782
transform 1 0 13632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_143
timestamp 1679581782
transform 1 0 14304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_150
timestamp 1679581782
transform 1 0 14976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_157
timestamp 1679581782
transform 1 0 15648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_164
timestamp 1679581782
transform 1 0 16320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_171
timestamp 1679581782
transform 1 0 16992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_178
timestamp 1679581782
transform 1 0 17664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_185
timestamp 1679581782
transform 1 0 18336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_192
timestamp 1679581782
transform 1 0 19008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_199
timestamp 1679581782
transform 1 0 19680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_206
timestamp 1679581782
transform 1 0 20352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_213
timestamp 1679581782
transform 1 0 21024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_220
timestamp 1679581782
transform 1 0 21696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_227
timestamp 1679581782
transform 1 0 22368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_234
timestamp 1679581782
transform 1 0 23040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_241
timestamp 1679581782
transform 1 0 23712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_248
timestamp 1679581782
transform 1 0 24384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_255
timestamp 1679581782
transform 1 0 25056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_262
timestamp 1679581782
transform 1 0 25728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_269
timestamp 1679581782
transform 1 0 26400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_276
timestamp 1679581782
transform 1 0 27072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_283
timestamp 1679581782
transform 1 0 27744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_290
timestamp 1679581782
transform 1 0 28416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_297
timestamp 1679581782
transform 1 0 29088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_304
timestamp 1679581782
transform 1 0 29760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_311
timestamp 1679581782
transform 1 0 30432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_318
timestamp 1679581782
transform 1 0 31104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_325
timestamp 1679581782
transform 1 0 31776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_332
timestamp 1679581782
transform 1 0 32448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_339
timestamp 1679581782
transform 1 0 33120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_346
timestamp 1679581782
transform 1 0 33792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_353
timestamp 1679581782
transform 1 0 34464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_360
timestamp 1679581782
transform 1 0 35136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_367
timestamp 1679577901
transform 1 0 35808 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_371
timestamp 1677579658
transform 1 0 36192 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_430
timestamp 1677580104
transform 1 0 41856 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_436
timestamp 1679581782
transform 1 0 42432 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_443
timestamp 1677580104
transform 1 0 43104 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_459
timestamp 1679581782
transform 1 0 44640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_466
timestamp 1679581782
transform 1 0 45312 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_473
timestamp 1677580104
transform 1 0 45984 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_507
timestamp 1679577901
transform 1 0 49248 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_511
timestamp 1677580104
transform 1 0 49632 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_540
timestamp 1677579658
transform 1 0 52416 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_555
timestamp 1679577901
transform 1 0 53856 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_563
timestamp 1679581782
transform 1 0 54624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_570
timestamp 1679581782
transform 1 0 55296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_577
timestamp 1679581782
transform 1 0 55968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_584
timestamp 1679581782
transform 1 0 56640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_625
timestamp 1679581782
transform 1 0 60576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_632
timestamp 1679581782
transform 1 0 61248 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_639
timestamp 1677580104
transform 1 0 61920 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_645
timestamp 1679581782
transform 1 0 62496 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_652
timestamp 1677580104
transform 1 0 63168 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_659
timestamp 1677580104
transform 1 0 63840 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_661
timestamp 1677579658
transform 1 0 64032 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_672
timestamp 1677579658
transform 1 0 65088 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_724
timestamp 1677580104
transform 1 0 70080 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_726
timestamp 1677579658
transform 1 0 70272 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_754
timestamp 1679577901
transform 1 0 72960 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_785
timestamp 1677579658
transform 1 0 75936 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_4
timestamp 1677579658
transform 1 0 960 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_40
timestamp 1679577901
transform 1 0 4416 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_48
timestamp 1679581782
transform 1 0 5184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_55
timestamp 1679581782
transform 1 0 5856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_62
timestamp 1679581782
transform 1 0 6528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_69
timestamp 1679581782
transform 1 0 7200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_76
timestamp 1679581782
transform 1 0 7872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_83
timestamp 1679581782
transform 1 0 8544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_90
timestamp 1679581782
transform 1 0 9216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_97
timestamp 1679581782
transform 1 0 9888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_104
timestamp 1679581782
transform 1 0 10560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_111
timestamp 1679581782
transform 1 0 11232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_118
timestamp 1679581782
transform 1 0 11904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_125
timestamp 1679581782
transform 1 0 12576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_132
timestamp 1679581782
transform 1 0 13248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_139
timestamp 1679581782
transform 1 0 13920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_146
timestamp 1679581782
transform 1 0 14592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_153
timestamp 1679581782
transform 1 0 15264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_160
timestamp 1679581782
transform 1 0 15936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_167
timestamp 1679581782
transform 1 0 16608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_174
timestamp 1679581782
transform 1 0 17280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_181
timestamp 1679581782
transform 1 0 17952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_188
timestamp 1679581782
transform 1 0 18624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_195
timestamp 1679581782
transform 1 0 19296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_202
timestamp 1679581782
transform 1 0 19968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_209
timestamp 1679581782
transform 1 0 20640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_216
timestamp 1679581782
transform 1 0 21312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_223
timestamp 1679581782
transform 1 0 21984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_230
timestamp 1679581782
transform 1 0 22656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_237
timestamp 1679581782
transform 1 0 23328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_244
timestamp 1679581782
transform 1 0 24000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_251
timestamp 1679581782
transform 1 0 24672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_258
timestamp 1679581782
transform 1 0 25344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_265
timestamp 1679581782
transform 1 0 26016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_272
timestamp 1679581782
transform 1 0 26688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_279
timestamp 1679581782
transform 1 0 27360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_286
timestamp 1679581782
transform 1 0 28032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_293
timestamp 1679581782
transform 1 0 28704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_300
timestamp 1679581782
transform 1 0 29376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_307
timestamp 1679581782
transform 1 0 30048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_314
timestamp 1679581782
transform 1 0 30720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_321
timestamp 1679581782
transform 1 0 31392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_328
timestamp 1679581782
transform 1 0 32064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_335
timestamp 1679581782
transform 1 0 32736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_342
timestamp 1679581782
transform 1 0 33408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_349
timestamp 1679581782
transform 1 0 34080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_356
timestamp 1679581782
transform 1 0 34752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_363
timestamp 1679577901
transform 1 0 35424 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_367
timestamp 1677579658
transform 1 0 35808 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_407
timestamp 1677579658
transform 1 0 39648 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_412
timestamp 1679581782
transform 1 0 40128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_419
timestamp 1679577901
transform 1 0 40800 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_423
timestamp 1677580104
transform 1 0 41184 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_439
timestamp 1679577901
transform 1 0 42720 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_443
timestamp 1677579658
transform 1 0 43104 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_480
timestamp 1677580104
transform 1 0 46656 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_486
timestamp 1679577901
transform 1 0 47232 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_521
timestamp 1677579658
transform 1 0 50592 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_527
timestamp 1677579658
transform 1 0 51168 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_536
timestamp 1679581782
transform 1 0 52032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_543
timestamp 1679577901
transform 1 0 52704 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_547
timestamp 1677580104
transform 1 0 53088 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_618
timestamp 1679581782
transform 1 0 59904 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_625
timestamp 1677580104
transform 1 0 60576 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_627
timestamp 1677579658
transform 1 0 60768 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_655
timestamp 1679577901
transform 1 0 63456 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_663
timestamp 1677580104
transform 1 0 64224 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_665
timestamp 1677579658
transform 1 0 64416 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_675
timestamp 1679577901
transform 1 0 65376 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_683
timestamp 1679581782
transform 1 0 66144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_690
timestamp 1679581782
transform 1 0 66816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_697
timestamp 1679581782
transform 1 0 67488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_704
timestamp 1679577901
transform 1 0 68160 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_721
timestamp 1677579658
transform 1 0 69792 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_726
timestamp 1677580104
transform 1 0 70272 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_740
timestamp 1679581782
transform 1 0 71616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_747
timestamp 1679577901
transform 1 0 72288 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_751
timestamp 1677580104
transform 1 0 72672 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_757
timestamp 1679581782
transform 1 0 73248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_764
timestamp 1679581782
transform 1 0 73920 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_794
timestamp 1677580104
transform 1 0 76800 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_800
timestamp 1677580104
transform 1 0 77376 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_806
timestamp 1679581782
transform 1 0 77952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_813
timestamp 1679581782
transform 1 0 78624 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_820
timestamp 1677580104
transform 1 0 79296 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_822
timestamp 1677579658
transform 1 0 79488 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_4
timestamp 1677580104
transform 1 0 960 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_19
timestamp 1679581782
transform 1 0 2400 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_26
timestamp 1677579658
transform 1 0 3072 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_37
timestamp 1677580104
transform 1 0 4128 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_39
timestamp 1677579658
transform 1 0 4320 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_72
timestamp 1679581782
transform 1 0 7488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_79
timestamp 1679581782
transform 1 0 8160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_86
timestamp 1679581782
transform 1 0 8832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_93
timestamp 1679581782
transform 1 0 9504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_100
timestamp 1679581782
transform 1 0 10176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_107
timestamp 1679581782
transform 1 0 10848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_114
timestamp 1679581782
transform 1 0 11520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_121
timestamp 1679581782
transform 1 0 12192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_128
timestamp 1679581782
transform 1 0 12864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_135
timestamp 1679581782
transform 1 0 13536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_142
timestamp 1679581782
transform 1 0 14208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_149
timestamp 1679581782
transform 1 0 14880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_156
timestamp 1679581782
transform 1 0 15552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_163
timestamp 1679581782
transform 1 0 16224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_170
timestamp 1679581782
transform 1 0 16896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_177
timestamp 1679581782
transform 1 0 17568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_184
timestamp 1679581782
transform 1 0 18240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_191
timestamp 1679581782
transform 1 0 18912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_198
timestamp 1679581782
transform 1 0 19584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_205
timestamp 1679581782
transform 1 0 20256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_212
timestamp 1679581782
transform 1 0 20928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_219
timestamp 1679581782
transform 1 0 21600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_226
timestamp 1679581782
transform 1 0 22272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_233
timestamp 1679581782
transform 1 0 22944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_240
timestamp 1679581782
transform 1 0 23616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_247
timestamp 1679581782
transform 1 0 24288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_254
timestamp 1679581782
transform 1 0 24960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_261
timestamp 1679581782
transform 1 0 25632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_268
timestamp 1679581782
transform 1 0 26304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_275
timestamp 1679581782
transform 1 0 26976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_282
timestamp 1679581782
transform 1 0 27648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_289
timestamp 1679581782
transform 1 0 28320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_296
timestamp 1679581782
transform 1 0 28992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_303
timestamp 1679581782
transform 1 0 29664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_310
timestamp 1679581782
transform 1 0 30336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_317
timestamp 1679581782
transform 1 0 31008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_324
timestamp 1679581782
transform 1 0 31680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_331
timestamp 1679581782
transform 1 0 32352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_338
timestamp 1679581782
transform 1 0 33024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_345
timestamp 1679577901
transform 1 0 33696 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_349
timestamp 1677580104
transform 1 0 34080 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_355
timestamp 1677579658
transform 1 0 34656 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_366
timestamp 1677580104
transform 1 0 35712 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_368
timestamp 1677579658
transform 1 0 35904 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_379
timestamp 1679581782
transform 1 0 36960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_386
timestamp 1679577901
transform 1 0 37632 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_409
timestamp 1679581782
transform 1 0 39840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_416
timestamp 1679581782
transform 1 0 40512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_423
timestamp 1679577901
transform 1 0 41184 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_427
timestamp 1677580104
transform 1 0 41568 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_465
timestamp 1679581782
transform 1 0 45216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_486
timestamp 1679581782
transform 1 0 47232 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_493
timestamp 1677580104
transform 1 0 47904 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_495
timestamp 1677579658
transform 1 0 48096 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_501
timestamp 1679577901
transform 1 0 48672 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_514
timestamp 1677580104
transform 1 0 49920 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_536
timestamp 1679577901
transform 1 0 52032 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_544
timestamp 1679581782
transform 1 0 52800 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_551
timestamp 1677580104
transform 1 0 53472 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_557
timestamp 1679581782
transform 1 0 54048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_564
timestamp 1679577901
transform 1 0 54720 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_568
timestamp 1677580104
transform 1 0 55104 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_574
timestamp 1679577901
transform 1 0 55680 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_587
timestamp 1677580104
transform 1 0 56928 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_589
timestamp 1677579658
transform 1 0 57120 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_604
timestamp 1677580104
transform 1 0 58560 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_642
timestamp 1679577901
transform 1 0 62208 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_646
timestamp 1677579658
transform 1 0 62592 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_652
timestamp 1677579658
transform 1 0 63168 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_668
timestamp 1679577901
transform 1 0 64704 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_672
timestamp 1677580104
transform 1 0 65088 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_678
timestamp 1679581782
transform 1 0 65664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_685
timestamp 1679581782
transform 1 0 66336 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_692
timestamp 1677580104
transform 1 0 67008 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_694
timestamp 1677579658
transform 1 0 67200 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_699
timestamp 1679581782
transform 1 0 67680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_706
timestamp 1679577901
transform 1 0 68352 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_710
timestamp 1677579658
transform 1 0 68736 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_716
timestamp 1677579658
transform 1 0 69312 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_731
timestamp 1679581782
transform 1 0 70752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_738
timestamp 1679581782
transform 1 0 71424 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_745
timestamp 1677580104
transform 1 0 72096 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_747
timestamp 1677579658
transform 1 0 72288 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_775
timestamp 1677580104
transform 1 0 74976 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_787
timestamp 1677580104
transform 1 0 76128 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_798
timestamp 1677579658
transform 1 0 77184 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_803
timestamp 1679581782
transform 1 0 77664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_810
timestamp 1679581782
transform 1 0 78336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_817
timestamp 1679577901
transform 1 0 79008 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_821
timestamp 1677580104
transform 1 0 79392 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_4
timestamp 1677579658
transform 1 0 960 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_27
timestamp 1679581782
transform 1 0 3168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_34
timestamp 1679577901
transform 1 0 3840 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_38
timestamp 1677580104
transform 1 0 4224 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_59
timestamp 1679581782
transform 1 0 6240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_66
timestamp 1679581782
transform 1 0 6912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_73
timestamp 1679581782
transform 1 0 7584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_80
timestamp 1679581782
transform 1 0 8256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_87
timestamp 1679581782
transform 1 0 8928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_94
timestamp 1679581782
transform 1 0 9600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_101
timestamp 1679581782
transform 1 0 10272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_108
timestamp 1679581782
transform 1 0 10944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_115
timestamp 1679581782
transform 1 0 11616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_122
timestamp 1679581782
transform 1 0 12288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_129
timestamp 1679581782
transform 1 0 12960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_136
timestamp 1679581782
transform 1 0 13632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_143
timestamp 1679581782
transform 1 0 14304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_150
timestamp 1679581782
transform 1 0 14976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_157
timestamp 1679581782
transform 1 0 15648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_164
timestamp 1679581782
transform 1 0 16320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_171
timestamp 1679581782
transform 1 0 16992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_178
timestamp 1679581782
transform 1 0 17664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_185
timestamp 1679581782
transform 1 0 18336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_192
timestamp 1679581782
transform 1 0 19008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_199
timestamp 1679581782
transform 1 0 19680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_206
timestamp 1679581782
transform 1 0 20352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_213
timestamp 1679581782
transform 1 0 21024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_220
timestamp 1679581782
transform 1 0 21696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_227
timestamp 1679581782
transform 1 0 22368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_234
timestamp 1679581782
transform 1 0 23040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_241
timestamp 1679581782
transform 1 0 23712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_248
timestamp 1679581782
transform 1 0 24384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_255
timestamp 1679581782
transform 1 0 25056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_262
timestamp 1679581782
transform 1 0 25728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_269
timestamp 1679581782
transform 1 0 26400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_276
timestamp 1679581782
transform 1 0 27072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_283
timestamp 1679581782
transform 1 0 27744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_290
timestamp 1679581782
transform 1 0 28416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_297
timestamp 1679581782
transform 1 0 29088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_304
timestamp 1679581782
transform 1 0 29760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_311
timestamp 1679581782
transform 1 0 30432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_318
timestamp 1679581782
transform 1 0 31104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_325
timestamp 1679581782
transform 1 0 31776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_332
timestamp 1679581782
transform 1 0 32448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_339
timestamp 1679581782
transform 1 0 33120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_387
timestamp 1679581782
transform 1 0 37728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_394
timestamp 1679577901
transform 1 0 38400 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_398
timestamp 1677580104
transform 1 0 38784 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_427
timestamp 1679577901
transform 1 0 41568 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_431
timestamp 1677580104
transform 1 0 41952 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_437
timestamp 1677580104
transform 1 0 42528 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_443
timestamp 1679581782
transform 1 0 43104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_450
timestamp 1679581782
transform 1 0 43776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_457
timestamp 1679581782
transform 1 0 44448 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_464
timestamp 1677580104
transform 1 0 45120 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_466
timestamp 1677579658
transform 1 0 45312 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_517
timestamp 1679581782
transform 1 0 50208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_524
timestamp 1679581782
transform 1 0 50880 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_562
timestamp 1677580104
transform 1 0 54528 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_564
timestamp 1677579658
transform 1 0 54720 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_592
timestamp 1679577901
transform 1 0 57408 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_604
timestamp 1679581782
transform 1 0 58560 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_615
timestamp 1677579658
transform 1 0 59616 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_620
timestamp 1679581782
transform 1 0 60096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_627
timestamp 1679577901
transform 1 0 60768 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_631
timestamp 1677579658
transform 1 0 61152 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_637
timestamp 1677580104
transform 1 0 61728 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_639
timestamp 1677579658
transform 1 0 61920 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_645
timestamp 1679577901
transform 1 0 62496 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_649
timestamp 1677579658
transform 1 0 62880 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_655
timestamp 1679581782
transform 1 0 63456 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_662
timestamp 1677580104
transform 1 0 64128 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_754
timestamp 1679581782
transform 1 0 72960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_761
timestamp 1679577901
transform 1 0 73632 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_765
timestamp 1677580104
transform 1 0 74016 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_777
timestamp 1679581782
transform 1 0 75168 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_784
timestamp 1677579658
transform 1 0 75840 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_789
timestamp 1679577901
transform 1 0 76320 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_793
timestamp 1677579658
transform 1 0 76704 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_821
timestamp 1677580104
transform 1 0 79392 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_4
timestamp 1677580104
transform 1 0 960 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_42
timestamp 1677580104
transform 1 0 4608 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_44
timestamp 1677579658
transform 1 0 4800 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_66
timestamp 1679581782
transform 1 0 6912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_73
timestamp 1679581782
transform 1 0 7584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_80
timestamp 1679581782
transform 1 0 8256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_87
timestamp 1679581782
transform 1 0 8928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_94
timestamp 1679581782
transform 1 0 9600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_101
timestamp 1679581782
transform 1 0 10272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_108
timestamp 1679581782
transform 1 0 10944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_115
timestamp 1679581782
transform 1 0 11616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_122
timestamp 1679581782
transform 1 0 12288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_129
timestamp 1679581782
transform 1 0 12960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_136
timestamp 1679581782
transform 1 0 13632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_143
timestamp 1679581782
transform 1 0 14304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_150
timestamp 1679581782
transform 1 0 14976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_157
timestamp 1679581782
transform 1 0 15648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_164
timestamp 1679581782
transform 1 0 16320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_171
timestamp 1679581782
transform 1 0 16992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_178
timestamp 1679581782
transform 1 0 17664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_185
timestamp 1679581782
transform 1 0 18336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_192
timestamp 1679581782
transform 1 0 19008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_199
timestamp 1679581782
transform 1 0 19680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_206
timestamp 1679581782
transform 1 0 20352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_213
timestamp 1679581782
transform 1 0 21024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_220
timestamp 1679581782
transform 1 0 21696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_227
timestamp 1679581782
transform 1 0 22368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_234
timestamp 1679581782
transform 1 0 23040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_241
timestamp 1679581782
transform 1 0 23712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_248
timestamp 1679581782
transform 1 0 24384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_255
timestamp 1679581782
transform 1 0 25056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_262
timestamp 1679581782
transform 1 0 25728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_269
timestamp 1679581782
transform 1 0 26400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_276
timestamp 1679581782
transform 1 0 27072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_283
timestamp 1679581782
transform 1 0 27744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_290
timestamp 1679581782
transform 1 0 28416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_297
timestamp 1679581782
transform 1 0 29088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_304
timestamp 1679581782
transform 1 0 29760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_311
timestamp 1679581782
transform 1 0 30432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_318
timestamp 1679581782
transform 1 0 31104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_325
timestamp 1679577901
transform 1 0 31776 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_329
timestamp 1677579658
transform 1 0 32160 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_339
timestamp 1679581782
transform 1 0 33120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_346
timestamp 1679581782
transform 1 0 33792 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_353
timestamp 1677580104
transform 1 0 34464 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_355
timestamp 1677579658
transform 1 0 34656 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_361
timestamp 1679581782
transform 1 0 35232 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_368
timestamp 1677580104
transform 1 0 35904 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_409
timestamp 1679581782
transform 1 0 39840 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_416
timestamp 1677580104
transform 1 0 40512 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_422
timestamp 1679577901
transform 1 0 41088 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_431
timestamp 1679581782
transform 1 0 41952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_469
timestamp 1679577901
transform 1 0 45600 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_491
timestamp 1677579658
transform 1 0 47712 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_497
timestamp 1677580104
transform 1 0 48288 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_499
timestamp 1677579658
transform 1 0 48480 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_504
timestamp 1679577901
transform 1 0 48960 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_535
timestamp 1679581782
transform 1 0 51936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_542
timestamp 1679581782
transform 1 0 52608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_549
timestamp 1679581782
transform 1 0 53280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_556
timestamp 1679577901
transform 1 0 53952 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_565
timestamp 1677580104
transform 1 0 54816 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_572
timestamp 1679577901
transform 1 0 55488 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_576
timestamp 1677579658
transform 1 0 55872 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_587
timestamp 1679581782
transform 1 0 56928 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_594
timestamp 1677579658
transform 1 0 57600 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_610
timestamp 1679581782
transform 1 0 59136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_617
timestamp 1679581782
transform 1 0 59808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_624
timestamp 1679577901
transform 1 0 60480 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_628
timestamp 1677579658
transform 1 0 60864 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_648
timestamp 1679581782
transform 1 0 62784 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_655
timestamp 1677580104
transform 1 0 63456 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_657
timestamp 1677579658
transform 1 0 63648 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_668
timestamp 1679577901
transform 1 0 64704 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_676
timestamp 1679581782
transform 1 0 65472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_683
timestamp 1679581782
transform 1 0 66144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_690
timestamp 1679581782
transform 1 0 66816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_697
timestamp 1679581782
transform 1 0 67488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_704
timestamp 1679577901
transform 1 0 68160 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_718
timestamp 1677579658
transform 1 0 69504 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_727
timestamp 1679577901
transform 1 0 70368 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_731
timestamp 1677580104
transform 1 0 70752 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_737
timestamp 1679577901
transform 1 0 71328 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_777
timestamp 1677579658
transform 1 0 75168 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_788
timestamp 1677580104
transform 1 0 76224 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_799
timestamp 1677579658
transform 1 0 77280 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_804
timestamp 1679581782
transform 1 0 77760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679581782
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_818
timestamp 1679577901
transform 1 0 79104 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_822
timestamp 1677579658
transform 1 0 79488 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_0
timestamp 1679577901
transform 1 0 576 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_4
timestamp 1677579658
transform 1 0 960 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_13
timestamp 1679577901
transform 1 0 1824 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_17
timestamp 1677579658
transform 1 0 2208 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_27
timestamp 1679581782
transform 1 0 3168 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_44
timestamp 1677580104
transform 1 0 4800 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_73
timestamp 1679581782
transform 1 0 7584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_80
timestamp 1679581782
transform 1 0 8256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_87
timestamp 1679581782
transform 1 0 8928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_94
timestamp 1679581782
transform 1 0 9600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_101
timestamp 1679581782
transform 1 0 10272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_108
timestamp 1679581782
transform 1 0 10944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_115
timestamp 1679581782
transform 1 0 11616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_122
timestamp 1679581782
transform 1 0 12288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_129
timestamp 1679581782
transform 1 0 12960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_136
timestamp 1679581782
transform 1 0 13632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_143
timestamp 1679581782
transform 1 0 14304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_150
timestamp 1679581782
transform 1 0 14976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_157
timestamp 1679581782
transform 1 0 15648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_164
timestamp 1679581782
transform 1 0 16320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_171
timestamp 1679581782
transform 1 0 16992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_178
timestamp 1679581782
transform 1 0 17664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_185
timestamp 1679581782
transform 1 0 18336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_192
timestamp 1679581782
transform 1 0 19008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_199
timestamp 1679581782
transform 1 0 19680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_206
timestamp 1679581782
transform 1 0 20352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_213
timestamp 1679581782
transform 1 0 21024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_220
timestamp 1679581782
transform 1 0 21696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_227
timestamp 1679581782
transform 1 0 22368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_234
timestamp 1679581782
transform 1 0 23040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_241
timestamp 1679581782
transform 1 0 23712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_248
timestamp 1679581782
transform 1 0 24384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_255
timestamp 1679581782
transform 1 0 25056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_262
timestamp 1679581782
transform 1 0 25728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_269
timestamp 1679581782
transform 1 0 26400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_276
timestamp 1679581782
transform 1 0 27072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_283
timestamp 1679581782
transform 1 0 27744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_290
timestamp 1679581782
transform 1 0 28416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_297
timestamp 1679581782
transform 1 0 29088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_304
timestamp 1679577901
transform 1 0 29760 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_308
timestamp 1677580104
transform 1 0 30144 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_314
timestamp 1679581782
transform 1 0 30720 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_326
timestamp 1677579658
transform 1 0 31872 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_364
timestamp 1679581782
transform 1 0 35520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679581782
transform 1 0 36192 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_378
timestamp 1677579658
transform 1 0 36864 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_397
timestamp 1679577901
transform 1 0 38688 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_406
timestamp 1677580104
transform 1 0 39552 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_454
timestamp 1679577901
transform 1 0 44160 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_17_485
timestamp 1679577901
transform 1 0 47136 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_494
timestamp 1679581782
transform 1 0 48000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_501
timestamp 1679581782
transform 1 0 48672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_508
timestamp 1679581782
transform 1 0 49344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_515
timestamp 1679581782
transform 1 0 50016 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_548
timestamp 1677579658
transform 1 0 53184 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_585
timestamp 1679581782
transform 1 0 56736 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_592
timestamp 1677580104
transform 1 0 57408 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_594
timestamp 1677579658
transform 1 0 57600 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_626
timestamp 1677579658
transform 1 0 60672 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_663
timestamp 1679577901
transform 1 0 64224 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_699
timestamp 1677580104
transform 1 0 67680 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_701
timestamp 1677579658
transform 1 0 67872 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_716
timestamp 1677580104
transform 1 0 69312 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_736
timestamp 1679581782
transform 1 0 71232 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_743
timestamp 1677580104
transform 1 0 71904 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_777
timestamp 1679577901
transform 1 0 75168 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_781
timestamp 1677580104
transform 1 0 75552 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_787
timestamp 1679581782
transform 1 0 76128 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_794
timestamp 1677579658
transform 1 0 76800 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_822
timestamp 1677579658
transform 1 0 79488 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_8
timestamp 1677579658
transform 1 0 1344 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_29
timestamp 1679581782
transform 1 0 3360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_36
timestamp 1679581782
transform 1 0 4032 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_43
timestamp 1677580104
transform 1 0 4704 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_45
timestamp 1677579658
transform 1 0 4896 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_50
timestamp 1679581782
transform 1 0 5376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_57
timestamp 1679581782
transform 1 0 6048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_64
timestamp 1679581782
transform 1 0 6720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_71
timestamp 1679581782
transform 1 0 7392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_78
timestamp 1679581782
transform 1 0 8064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_85
timestamp 1679581782
transform 1 0 8736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_92
timestamp 1679581782
transform 1 0 9408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_99
timestamp 1679581782
transform 1 0 10080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_106
timestamp 1679581782
transform 1 0 10752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_113
timestamp 1679581782
transform 1 0 11424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_120
timestamp 1679581782
transform 1 0 12096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_127
timestamp 1679581782
transform 1 0 12768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_134
timestamp 1679581782
transform 1 0 13440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_141
timestamp 1679581782
transform 1 0 14112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_148
timestamp 1679581782
transform 1 0 14784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_155
timestamp 1679581782
transform 1 0 15456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_162
timestamp 1679581782
transform 1 0 16128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_169
timestamp 1679581782
transform 1 0 16800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_176
timestamp 1679581782
transform 1 0 17472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_183
timestamp 1679581782
transform 1 0 18144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_190
timestamp 1679581782
transform 1 0 18816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_197
timestamp 1679581782
transform 1 0 19488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_204
timestamp 1679581782
transform 1 0 20160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_211
timestamp 1679581782
transform 1 0 20832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_218
timestamp 1679581782
transform 1 0 21504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_225
timestamp 1679581782
transform 1 0 22176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_232
timestamp 1679581782
transform 1 0 22848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_239
timestamp 1679581782
transform 1 0 23520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_246
timestamp 1679581782
transform 1 0 24192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_253
timestamp 1679581782
transform 1 0 24864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_260
timestamp 1679581782
transform 1 0 25536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_267
timestamp 1679581782
transform 1 0 26208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_274
timestamp 1679581782
transform 1 0 26880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_281
timestamp 1679581782
transform 1 0 27552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_288
timestamp 1679581782
transform 1 0 28224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_295
timestamp 1679581782
transform 1 0 28896 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_302
timestamp 1677580104
transform 1 0 29568 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_304
timestamp 1677579658
transform 1 0 29760 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_332
timestamp 1677580104
transform 1 0 32448 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_339
timestamp 1677580104
transform 1 0 33120 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_341
timestamp 1677579658
transform 1 0 33312 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_346
timestamp 1679581782
transform 1 0 33792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_353
timestamp 1679581782
transform 1 0 34464 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_360
timestamp 1677580104
transform 1 0 35136 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_366
timestamp 1677580104
transform 1 0 35712 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_415
timestamp 1679581782
transform 1 0 40416 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_422
timestamp 1677579658
transform 1 0 41088 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_428
timestamp 1679581782
transform 1 0 41664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_435
timestamp 1679577901
transform 1 0 42336 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_448
timestamp 1679581782
transform 1 0 43584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_455
timestamp 1679581782
transform 1 0 44256 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_462
timestamp 1677579658
transform 1 0 44928 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_467
timestamp 1677579658
transform 1 0 45408 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_486
timestamp 1677579658
transform 1 0 47232 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_491
timestamp 1677580104
transform 1 0 47712 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_520
timestamp 1677580104
transform 1 0 50496 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_549
timestamp 1679581782
transform 1 0 53280 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_556
timestamp 1677580104
transform 1 0 53952 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_558
timestamp 1677579658
transform 1 0 54144 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_563
timestamp 1679581782
transform 1 0 54624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_570
timestamp 1679577901
transform 1 0 55296 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_574
timestamp 1677580104
transform 1 0 55680 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_595
timestamp 1679581782
transform 1 0 57696 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_602
timestamp 1677580104
transform 1 0 58368 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_608
timestamp 1679581782
transform 1 0 58944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_615
timestamp 1679581782
transform 1 0 59616 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_622
timestamp 1677580104
transform 1 0 60288 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_649
timestamp 1679581782
transform 1 0 62880 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_656
timestamp 1677579658
transform 1 0 63552 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_676
timestamp 1679577901
transform 1 0 65472 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_684
timestamp 1679581782
transform 1 0 66240 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_691
timestamp 1677580104
transform 1 0 66912 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_724
timestamp 1677580104
transform 1 0 70080 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_753
timestamp 1679581782
transform 1 0 72864 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_780
timestamp 1677579658
transform 1 0 75456 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_786
timestamp 1677579658
transform 1 0 76032 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_821
timestamp 1677580104
transform 1 0 79392 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_35
timestamp 1677580104
transform 1 0 3936 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_50
timestamp 1679581782
transform 1 0 5376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_57
timestamp 1679581782
transform 1 0 6048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_64
timestamp 1679581782
transform 1 0 6720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_71
timestamp 1679581782
transform 1 0 7392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_78
timestamp 1679581782
transform 1 0 8064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_85
timestamp 1679581782
transform 1 0 8736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_92
timestamp 1679581782
transform 1 0 9408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_99
timestamp 1679581782
transform 1 0 10080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_106
timestamp 1679581782
transform 1 0 10752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_113
timestamp 1679581782
transform 1 0 11424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_120
timestamp 1679581782
transform 1 0 12096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_127
timestamp 1679581782
transform 1 0 12768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_134
timestamp 1679581782
transform 1 0 13440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_141
timestamp 1679581782
transform 1 0 14112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_148
timestamp 1679581782
transform 1 0 14784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_155
timestamp 1679581782
transform 1 0 15456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_162
timestamp 1679581782
transform 1 0 16128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_169
timestamp 1679581782
transform 1 0 16800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_176
timestamp 1679581782
transform 1 0 17472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_183
timestamp 1679581782
transform 1 0 18144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_190
timestamp 1679581782
transform 1 0 18816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_197
timestamp 1679581782
transform 1 0 19488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_204
timestamp 1679581782
transform 1 0 20160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_211
timestamp 1679581782
transform 1 0 20832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_218
timestamp 1679581782
transform 1 0 21504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_225
timestamp 1679581782
transform 1 0 22176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_232
timestamp 1679581782
transform 1 0 22848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_239
timestamp 1679581782
transform 1 0 23520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_246
timestamp 1679581782
transform 1 0 24192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_253
timestamp 1679581782
transform 1 0 24864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_260
timestamp 1679581782
transform 1 0 25536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_267
timestamp 1679581782
transform 1 0 26208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_274
timestamp 1679581782
transform 1 0 26880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_281
timestamp 1679581782
transform 1 0 27552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_288
timestamp 1679581782
transform 1 0 28224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_295
timestamp 1679581782
transform 1 0 28896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_302
timestamp 1679581782
transform 1 0 29568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_309
timestamp 1679581782
transform 1 0 30240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_316
timestamp 1679577901
transform 1 0 30912 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_320
timestamp 1677579658
transform 1 0 31296 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_325
timestamp 1677579658
transform 1 0 31776 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_330
timestamp 1679577901
transform 1 0 32256 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_334
timestamp 1677579658
transform 1 0 32640 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_350
timestamp 1677580104
transform 1 0 34176 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_393
timestamp 1679581782
transform 1 0 38304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_423
timestamp 1679577901
transform 1 0 41184 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_427
timestamp 1677580104
transform 1 0 41568 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_434
timestamp 1679581782
transform 1 0 42240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679581782
transform 1 0 42912 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_448
timestamp 1677579658
transform 1 0 43584 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_453
timestamp 1679581782
transform 1 0 44064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_460
timestamp 1679577901
transform 1 0 44736 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_464
timestamp 1677580104
transform 1 0 45120 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_480
timestamp 1677579658
transform 1 0 46656 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_495
timestamp 1677580104
transform 1 0 48096 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_497
timestamp 1677579658
transform 1 0 48288 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_502
timestamp 1677580104
transform 1 0 48768 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_504
timestamp 1677579658
transform 1 0 48960 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_509
timestamp 1677580104
transform 1 0 49440 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_516
timestamp 1679581782
transform 1 0 50112 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_528
timestamp 1677580104
transform 1 0 51264 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_535
timestamp 1677579658
transform 1 0 51936 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_546
timestamp 1677579658
transform 1 0 52992 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_574
timestamp 1679581782
transform 1 0 55680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_581
timestamp 1679581782
transform 1 0 56352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_615
timestamp 1679581782
transform 1 0 59616 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_622
timestamp 1677580104
transform 1 0 60288 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679581782
transform 1 0 63072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679581782
transform 1 0 63744 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_665
timestamp 1677580104
transform 1 0 64416 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_667
timestamp 1677579658
transform 1 0 64608 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_672
timestamp 1677580104
transform 1 0 65088 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_674
timestamp 1677579658
transform 1 0 65280 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_706
timestamp 1677580104
transform 1 0 68352 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_708
timestamp 1677579658
transform 1 0 68544 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_713
timestamp 1679577901
transform 1 0 69024 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_717
timestamp 1677580104
transform 1 0 69408 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_740
timestamp 1679581782
transform 1 0 71616 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_747
timestamp 1677580104
transform 1 0 72288 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_749
timestamp 1677579658
transform 1 0 72480 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_754
timestamp 1679581782
transform 1 0 72960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_761
timestamp 1679581782
transform 1 0 73632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_768
timestamp 1679581782
transform 1 0 74304 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_775
timestamp 1677579658
transform 1 0 74976 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_780
timestamp 1679581782
transform 1 0 75456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_787
timestamp 1679577901
transform 1 0 76128 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_791
timestamp 1677579658
transform 1 0 76512 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_796
timestamp 1679581782
transform 1 0 76992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_803
timestamp 1679581782
transform 1 0 77664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_810
timestamp 1679581782
transform 1 0 78336 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_817
timestamp 1677580104
transform 1 0 79008 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_819
timestamp 1677579658
transform 1 0 79200 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_4
timestamp 1679577901
transform 1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_8
timestamp 1677579658
transform 1 0 1344 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_13
timestamp 1677579658
transform 1 0 1824 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_26
timestamp 1677580104
transform 1 0 3072 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_32
timestamp 1679577901
transform 1 0 3648 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_36
timestamp 1677579658
transform 1 0 4032 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_68
timestamp 1679581782
transform 1 0 7104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_75
timestamp 1679581782
transform 1 0 7776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_82
timestamp 1679581782
transform 1 0 8448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_89
timestamp 1679581782
transform 1 0 9120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_96
timestamp 1679581782
transform 1 0 9792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_103
timestamp 1679581782
transform 1 0 10464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_110
timestamp 1679581782
transform 1 0 11136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_117
timestamp 1679581782
transform 1 0 11808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_124
timestamp 1679581782
transform 1 0 12480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_131
timestamp 1679581782
transform 1 0 13152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_138
timestamp 1679581782
transform 1 0 13824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_145
timestamp 1679581782
transform 1 0 14496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_152
timestamp 1679581782
transform 1 0 15168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_159
timestamp 1679581782
transform 1 0 15840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_166
timestamp 1679581782
transform 1 0 16512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_173
timestamp 1679581782
transform 1 0 17184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_180
timestamp 1679581782
transform 1 0 17856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_187
timestamp 1679581782
transform 1 0 18528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_194
timestamp 1679581782
transform 1 0 19200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_201
timestamp 1679581782
transform 1 0 19872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_208
timestamp 1679581782
transform 1 0 20544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_215
timestamp 1679581782
transform 1 0 21216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_222
timestamp 1679581782
transform 1 0 21888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_229
timestamp 1679581782
transform 1 0 22560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_236
timestamp 1679581782
transform 1 0 23232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_243
timestamp 1679581782
transform 1 0 23904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_250
timestamp 1679581782
transform 1 0 24576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_257
timestamp 1679581782
transform 1 0 25248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_264
timestamp 1679581782
transform 1 0 25920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_271
timestamp 1679581782
transform 1 0 26592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_282
timestamp 1679581782
transform 1 0 27648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_289
timestamp 1679581782
transform 1 0 28320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_296
timestamp 1679581782
transform 1 0 28992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_303
timestamp 1679581782
transform 1 0 29664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_310
timestamp 1679577901
transform 1 0 30336 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_314
timestamp 1677580104
transform 1 0 30720 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_357
timestamp 1679581782
transform 1 0 34848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_364
timestamp 1679581782
transform 1 0 35520 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_371
timestamp 1677579658
transform 1 0 36192 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_391
timestamp 1679581782
transform 1 0 38112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_398
timestamp 1679581782
transform 1 0 38784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_405
timestamp 1679577901
transform 1 0 39456 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_471
timestamp 1677579658
transform 1 0 45792 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_485
timestamp 1679581782
transform 1 0 47136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_492
timestamp 1679581782
transform 1 0 47808 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_499
timestamp 1677579658
transform 1 0 48480 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_535
timestamp 1679577901
transform 1 0 51936 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_539
timestamp 1677580104
transform 1 0 52320 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_550
timestamp 1677580104
transform 1 0 53376 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_556
timestamp 1679577901
transform 1 0 53952 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_563
timestamp 1677579658
transform 1 0 54624 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_567
timestamp 1677580104
transform 1 0 55008 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_572
timestamp 1677579658
transform 1 0 55488 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_576
timestamp 1677580104
transform 1 0 55872 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_581
timestamp 1677579658
transform 1 0 56352 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_585
timestamp 1677579658
transform 1 0 56736 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_589
timestamp 1677579658
transform 1 0 57120 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_606
timestamp 1677579658
transform 1 0 58752 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_610
timestamp 1677579658
transform 1 0 59136 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_614
timestamp 1677579658
transform 1 0 59520 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_618
timestamp 1677579658
transform 1 0 59904 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_622
timestamp 1677580104
transform 1 0 60288 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_627
timestamp 1677580104
transform 1 0 60768 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_664
timestamp 1677579658
transform 1 0 64320 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_668
timestamp 1677580104
transform 1 0 64704 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_673
timestamp 1677579658
transform 1 0 65184 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_677
timestamp 1677579658
transform 1 0 65568 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_681
timestamp 1677579658
transform 1 0 65952 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_685
timestamp 1677579658
transform 1 0 66336 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_689
timestamp 1677580104
transform 1 0 66720 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_694
timestamp 1677579658
transform 1 0 67200 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_698
timestamp 1677579658
transform 1 0 67584 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_702
timestamp 1677579658
transform 1 0 67968 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_706
timestamp 1677579658
transform 1 0 68352 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_710
timestamp 1677580104
transform 1 0 68736 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_715
timestamp 1677579658
transform 1 0 69216 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_719
timestamp 1677579658
transform 1 0 69600 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_723
timestamp 1677579658
transform 1 0 69984 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_727
timestamp 1677579658
transform 1 0 70368 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_731
timestamp 1677579658
transform 1 0 70752 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_735
timestamp 1677579658
transform 1 0 71136 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_739
timestamp 1677580104
transform 1 0 71520 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_744
timestamp 1677579658
transform 1 0 72000 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_748
timestamp 1677579658
transform 1 0 72384 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_752
timestamp 1677579658
transform 1 0 72768 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_756
timestamp 1677579658
transform 1 0 73152 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_760
timestamp 1677579658
transform 1 0 73536 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_764
timestamp 1677580104
transform 1 0 73920 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_769
timestamp 1677579658
transform 1 0 74400 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_773
timestamp 1677579658
transform 1 0 74784 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_777
timestamp 1677579658
transform 1 0 75168 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_781
timestamp 1677579658
transform 1 0 75552 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_785
timestamp 1679577901
transform 1 0 75936 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_789
timestamp 1677579658
transform 1 0 76320 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_793
timestamp 1677579658
transform 1 0 76704 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_803
timestamp 1677579658
transform 1 0 77664 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_807
timestamp 1677579658
transform 1 0 78048 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_811
timestamp 1677579658
transform 1 0 78432 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_821
timestamp 1677580104
transform 1 0 79392 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_18
timestamp 1677579658
transform 1 0 2304 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_23
timestamp 1679581782
transform 1 0 2784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_30
timestamp 1679581782
transform 1 0 3456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_37
timestamp 1679581782
transform 1 0 4128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_44
timestamp 1679581782
transform 1 0 4800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_51
timestamp 1679581782
transform 1 0 5472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_58
timestamp 1679581782
transform 1 0 6144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_65
timestamp 1679581782
transform 1 0 6816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_72
timestamp 1679581782
transform 1 0 7488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_79
timestamp 1679581782
transform 1 0 8160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_86
timestamp 1679581782
transform 1 0 8832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_93
timestamp 1679581782
transform 1 0 9504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_100
timestamp 1679581782
transform 1 0 10176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_107
timestamp 1679581782
transform 1 0 10848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_114
timestamp 1679581782
transform 1 0 11520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_121
timestamp 1679581782
transform 1 0 12192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_128
timestamp 1679581782
transform 1 0 12864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_135
timestamp 1679581782
transform 1 0 13536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_142
timestamp 1679581782
transform 1 0 14208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_149
timestamp 1679581782
transform 1 0 14880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_156
timestamp 1679581782
transform 1 0 15552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_163
timestamp 1679581782
transform 1 0 16224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_170
timestamp 1679581782
transform 1 0 16896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_177
timestamp 1679581782
transform 1 0 17568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_184
timestamp 1679581782
transform 1 0 18240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_191
timestamp 1679581782
transform 1 0 18912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_198
timestamp 1679581782
transform 1 0 19584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_205
timestamp 1679581782
transform 1 0 20256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_212
timestamp 1679581782
transform 1 0 20928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_219
timestamp 1679581782
transform 1 0 21600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_226
timestamp 1679577901
transform 1 0 22272 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_238
timestamp 1677580104
transform 1 0 23424 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_244
timestamp 1679581782
transform 1 0 24000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_251
timestamp 1679581782
transform 1 0 24672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_258
timestamp 1679581782
transform 1 0 25344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_265
timestamp 1679581782
transform 1 0 26016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_304
timestamp 1679581782
transform 1 0 29760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_319
timestamp 1679581782
transform 1 0 31200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_326
timestamp 1679581782
transform 1 0 31872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_333
timestamp 1679581782
transform 1 0 32544 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_340
timestamp 1677579658
transform 1 0 33216 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_377
timestamp 1677579658
transform 1 0 36768 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_409
timestamp 1679581782
transform 1 0 39840 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_416
timestamp 1677580104
transform 1 0 40512 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_418
timestamp 1677579658
transform 1 0 40704 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_446
timestamp 1677580104
transform 1 0 43392 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_456
timestamp 1677579658
transform 1 0 44352 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_502
timestamp 1677580104
transform 1 0 48768 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_504
timestamp 1677579658
transform 1 0 48960 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_510
timestamp 1677580104
transform 1 0 49536 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_512
timestamp 1677579658
transform 1 0 49728 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_535
timestamp 1677580104
transform 1 0 51936 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_537
timestamp 1677579658
transform 1 0 52128 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_4
timestamp 1679577901
transform 1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_8
timestamp 1677579658
transform 1 0 1344 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_13
timestamp 1679581782
transform 1 0 1824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_20
timestamp 1679581782
transform 1 0 2496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_27
timestamp 1679581782
transform 1 0 3168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_34
timestamp 1679581782
transform 1 0 3840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_41
timestamp 1679581782
transform 1 0 4512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_48
timestamp 1679581782
transform 1 0 5184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_55
timestamp 1679581782
transform 1 0 5856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_62
timestamp 1679581782
transform 1 0 6528 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_69
timestamp 1677580104
transform 1 0 7200 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_71
timestamp 1677579658
transform 1 0 7392 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_86
timestamp 1679581782
transform 1 0 8832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_93
timestamp 1679581782
transform 1 0 9504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_100
timestamp 1679581782
transform 1 0 10176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_107
timestamp 1679581782
transform 1 0 10848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_114
timestamp 1679581782
transform 1 0 11520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_121
timestamp 1679581782
transform 1 0 12192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_128
timestamp 1679581782
transform 1 0 12864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_135
timestamp 1679581782
transform 1 0 13536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_142
timestamp 1679581782
transform 1 0 14208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_149
timestamp 1679581782
transform 1 0 14880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_156
timestamp 1679581782
transform 1 0 15552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_163
timestamp 1679581782
transform 1 0 16224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_170
timestamp 1679581782
transform 1 0 16896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_177
timestamp 1679581782
transform 1 0 17568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_184
timestamp 1679581782
transform 1 0 18240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_191
timestamp 1679581782
transform 1 0 18912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_198
timestamp 1679581782
transform 1 0 19584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_205
timestamp 1679581782
transform 1 0 20256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_212
timestamp 1679581782
transform 1 0 20928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_219
timestamp 1679577901
transform 1 0 21600 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_223
timestamp 1677580104
transform 1 0 21984 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_261
timestamp 1679581782
transform 1 0 25632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_286
timestamp 1679581782
transform 1 0 28032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_293
timestamp 1679581782
transform 1 0 28704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_300
timestamp 1679577901
transform 1 0 29376 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_304
timestamp 1677579658
transform 1 0 29760 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_337
timestamp 1677580104
transform 1 0 32928 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_339
timestamp 1677579658
transform 1 0 33120 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_344
timestamp 1679577901
transform 1 0 33600 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_348
timestamp 1677579658
transform 1 0 33984 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_353
timestamp 1677580104
transform 1 0 34464 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_359
timestamp 1679581782
transform 1 0 35040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_366
timestamp 1679577901
transform 1 0 35712 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_370
timestamp 1677580104
transform 1 0 36096 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_380
timestamp 1679581782
transform 1 0 37056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_391
timestamp 1679581782
transform 1 0 38112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_398
timestamp 1679581782
transform 1 0 38784 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_405
timestamp 1677580104
transform 1 0 39456 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_407
timestamp 1677579658
transform 1 0 39648 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_435
timestamp 1677580104
transform 1 0 42336 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_437
timestamp 1677579658
transform 1 0 42528 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_470
timestamp 1677580104
transform 1 0 45696 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_472
timestamp 1677579658
transform 1 0 45888 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_482
timestamp 1679581782
transform 1 0 46848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_489
timestamp 1679581782
transform 1 0 47520 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_505
timestamp 1677580104
transform 1 0 49056 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_507
timestamp 1677579658
transform 1 0 49248 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679581782
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679581782
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679581782
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679581782
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679581782
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_53
timestamp 1677580104
transform 1 0 5664 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_99
timestamp 1679581782
transform 1 0 10080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_106
timestamp 1679581782
transform 1 0 10752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_113
timestamp 1679581782
transform 1 0 11424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_120
timestamp 1679581782
transform 1 0 12096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_127
timestamp 1679581782
transform 1 0 12768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_134
timestamp 1679581782
transform 1 0 13440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_141
timestamp 1679581782
transform 1 0 14112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_148
timestamp 1679581782
transform 1 0 14784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_155
timestamp 1679581782
transform 1 0 15456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_162
timestamp 1679581782
transform 1 0 16128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_169
timestamp 1679581782
transform 1 0 16800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_176
timestamp 1679581782
transform 1 0 17472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_183
timestamp 1679581782
transform 1 0 18144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_190
timestamp 1679581782
transform 1 0 18816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_197
timestamp 1679581782
transform 1 0 19488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_204
timestamp 1679581782
transform 1 0 20160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_211
timestamp 1679577901
transform 1 0 20832 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_215
timestamp 1677580104
transform 1 0 21216 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_251
timestamp 1679577901
transform 1 0 24672 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_255
timestamp 1677580104
transform 1 0 25056 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_262
timestamp 1677579658
transform 1 0 25728 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_273
timestamp 1679581782
transform 1 0 26784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_280
timestamp 1679581782
transform 1 0 27456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_287
timestamp 1679577901
transform 1 0 28128 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_291
timestamp 1677579658
transform 1 0 28512 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_321
timestamp 1679577901
transform 1 0 31392 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_330
timestamp 1677580104
transform 1 0 32256 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_364
timestamp 1677579658
transform 1 0 35520 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_424
timestamp 1677580104
transform 1 0 41280 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_444
timestamp 1677580104
transform 1 0 43200 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_446
timestamp 1677579658
transform 1 0 43392 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_460
timestamp 1679581782
transform 1 0 44736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_467
timestamp 1679581782
transform 1 0 45408 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_478
timestamp 1677580104
transform 1 0 46464 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_485
timestamp 1677580104
transform 1 0 47136 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_492
timestamp 1677579658
transform 1 0 47808 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_511
timestamp 1677580104
transform 1 0 49632 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_517
timestamp 1677579658
transform 1 0 50208 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_530
timestamp 1679581782
transform 1 0 51456 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_537
timestamp 1677579658
transform 1 0 52128 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_64
timestamp 1679581782
transform 1 0 6720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_71
timestamp 1679581782
transform 1 0 7392 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_78
timestamp 1677580104
transform 1 0 8064 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_117
timestamp 1679581782
transform 1 0 11808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_124
timestamp 1679581782
transform 1 0 12480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_131
timestamp 1679581782
transform 1 0 13152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_138
timestamp 1679581782
transform 1 0 13824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_145
timestamp 1679581782
transform 1 0 14496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_152
timestamp 1679581782
transform 1 0 15168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_159
timestamp 1679581782
transform 1 0 15840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_166
timestamp 1679581782
transform 1 0 16512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_173
timestamp 1679581782
transform 1 0 17184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_180
timestamp 1679581782
transform 1 0 17856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_187
timestamp 1679581782
transform 1 0 18528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_194
timestamp 1679581782
transform 1 0 19200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_201
timestamp 1679581782
transform 1 0 19872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_208
timestamp 1679581782
transform 1 0 20544 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_215
timestamp 1677580104
transform 1 0 21216 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_217
timestamp 1677579658
transform 1 0 21408 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_258
timestamp 1677580104
transform 1 0 25344 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_260
timestamp 1677579658
transform 1 0 25536 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_292
timestamp 1679577901
transform 1 0 28608 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_296
timestamp 1677580104
transform 1 0 28992 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_325
timestamp 1677580104
transform 1 0 31776 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_327
timestamp 1677579658
transform 1 0 31968 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_333
timestamp 1677580104
transform 1 0 32544 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_335
timestamp 1677579658
transform 1 0 32736 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_350
timestamp 1679581782
transform 1 0 34176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_357
timestamp 1679581782
transform 1 0 34848 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_364
timestamp 1677579658
transform 1 0 35520 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_383
timestamp 1679581782
transform 1 0 37344 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_390
timestamp 1677579658
transform 1 0 38016 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_410
timestamp 1677580104
transform 1 0 39936 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_412
timestamp 1677579658
transform 1 0 40128 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_438
timestamp 1677579658
transform 1 0 42624 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_503
timestamp 1677579658
transform 1 0 48864 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_509
timestamp 1677579658
transform 1 0 49440 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_537
timestamp 1679581782
transform 1 0 52128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679581782
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679581782
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679581782
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679581782
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679581782
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679581782
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_81
timestamp 1679577901
transform 1 0 8352 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_85
timestamp 1677580104
transform 1 0 8736 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_91
timestamp 1679581782
transform 1 0 9312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_98
timestamp 1679581782
transform 1 0 9984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_105
timestamp 1679581782
transform 1 0 10656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_112
timestamp 1679581782
transform 1 0 11328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_119
timestamp 1679581782
transform 1 0 12000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_126
timestamp 1679581782
transform 1 0 12672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_133
timestamp 1679581782
transform 1 0 13344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_140
timestamp 1679581782
transform 1 0 14016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_147
timestamp 1679581782
transform 1 0 14688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_154
timestamp 1679581782
transform 1 0 15360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_161
timestamp 1679581782
transform 1 0 16032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_168
timestamp 1679581782
transform 1 0 16704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_175
timestamp 1679581782
transform 1 0 17376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_182
timestamp 1679581782
transform 1 0 18048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_189
timestamp 1679581782
transform 1 0 18720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_196
timestamp 1679581782
transform 1 0 19392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_203
timestamp 1679581782
transform 1 0 20064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_210
timestamp 1679581782
transform 1 0 20736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_217
timestamp 1679581782
transform 1 0 21408 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_224
timestamp 1677580104
transform 1 0 22080 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_235
timestamp 1677579658
transform 1 0 23136 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_240
timestamp 1679581782
transform 1 0 23616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_247
timestamp 1679581782
transform 1 0 24288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_254
timestamp 1679577901
transform 1 0 24960 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_262
timestamp 1679577901
transform 1 0 25728 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_266
timestamp 1677579658
transform 1 0 26112 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_280
timestamp 1677580104
transform 1 0 27456 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_282
timestamp 1677579658
transform 1 0 27648 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_297
timestamp 1679577901
transform 1 0 29088 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_301
timestamp 1677580104
transform 1 0 29472 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_307
timestamp 1679581782
transform 1 0 30048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_314
timestamp 1679577901
transform 1 0 30720 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_331
timestamp 1677580104
transform 1 0 32352 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_342
timestamp 1679581782
transform 1 0 33408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_349
timestamp 1679581782
transform 1 0 34080 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_356
timestamp 1677579658
transform 1 0 34752 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_362
timestamp 1677579658
transform 1 0 35328 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_373
timestamp 1679581782
transform 1 0 36384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_380
timestamp 1679577901
transform 1 0 37056 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_418
timestamp 1677580104
transform 1 0 40704 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_452
timestamp 1677580104
transform 1 0 43968 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_454
timestamp 1677579658
transform 1 0 44160 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_471
timestamp 1679581782
transform 1 0 45792 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_478
timestamp 1677580104
transform 1 0 46464 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_480
timestamp 1677579658
transform 1 0 46656 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_485
timestamp 1677579658
transform 1 0 47136 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_494
timestamp 1679581782
transform 1 0 48000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_501
timestamp 1679577901
transform 1 0 48672 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_509
timestamp 1679577901
transform 1 0 49440 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_513
timestamp 1677580104
transform 1 0 49824 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_519
timestamp 1679581782
transform 1 0 50400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_526
timestamp 1679581782
transform 1 0 51072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_533
timestamp 1679581782
transform 1 0 51744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_540
timestamp 1679577901
transform 1 0 52416 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679581782
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679581782
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679581782
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_46
timestamp 1679577901
transform 1 0 4992 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_53
timestamp 1679581782
transform 1 0 5664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679581782
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679581782
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679581782
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679581782
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679581782
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679581782
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679581782
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679581782
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679581782
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679581782
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679581782
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679581782
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679581782
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679581782
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679581782
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679581782
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679581782
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_256
timestamp 1679577901
transform 1 0 25152 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_260
timestamp 1677580104
transform 1 0 25536 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_289
timestamp 1677580104
transform 1 0 28320 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_291
timestamp 1677579658
transform 1 0 28512 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_297
timestamp 1677579658
transform 1 0 29088 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_329
timestamp 1677579658
transform 1 0 32160 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_357
timestamp 1679577901
transform 1 0 34848 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_361
timestamp 1677579658
transform 1 0 35232 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_389
timestamp 1677580104
transform 1 0 37920 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_391
timestamp 1677579658
transform 1 0 38112 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_424
timestamp 1677580104
transform 1 0 41280 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_435
timestamp 1679577901
transform 1 0 42336 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_439
timestamp 1677579658
transform 1 0 42720 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_452
timestamp 1677579658
transform 1 0 43968 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_457
timestamp 1677580104
transform 1 0 44448 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_459
timestamp 1677579658
transform 1 0 44640 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_465
timestamp 1677580104
transform 1 0 45216 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_481
timestamp 1679581782
transform 1 0 46752 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_488
timestamp 1677580104
transform 1 0 47424 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_34
timestamp 1679581782
transform 1 0 3840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_41
timestamp 1679581782
transform 1 0 4512 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_48
timestamp 1677580104
transform 1 0 5184 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_50
timestamp 1677579658
transform 1 0 5376 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_59
timestamp 1679581782
transform 1 0 6240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_66
timestamp 1679581782
transform 1 0 6912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_73
timestamp 1679581782
transform 1 0 7584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_80
timestamp 1679581782
transform 1 0 8256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_87
timestamp 1679581782
transform 1 0 8928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_94
timestamp 1679581782
transform 1 0 9600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_101
timestamp 1679581782
transform 1 0 10272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_108
timestamp 1679581782
transform 1 0 10944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_115
timestamp 1679581782
transform 1 0 11616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_122
timestamp 1679581782
transform 1 0 12288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_129
timestamp 1679581782
transform 1 0 12960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_136
timestamp 1679581782
transform 1 0 13632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_143
timestamp 1679581782
transform 1 0 14304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_150
timestamp 1679581782
transform 1 0 14976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_157
timestamp 1679581782
transform 1 0 15648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_164
timestamp 1679581782
transform 1 0 16320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_171
timestamp 1679581782
transform 1 0 16992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_178
timestamp 1679581782
transform 1 0 17664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_185
timestamp 1679581782
transform 1 0 18336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_192
timestamp 1679581782
transform 1 0 19008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_199
timestamp 1679581782
transform 1 0 19680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_206
timestamp 1679581782
transform 1 0 20352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_213
timestamp 1679581782
transform 1 0 21024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_220
timestamp 1679581782
transform 1 0 21696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_227
timestamp 1679581782
transform 1 0 22368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_234
timestamp 1679581782
transform 1 0 23040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_241
timestamp 1679581782
transform 1 0 23712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_248
timestamp 1679581782
transform 1 0 24384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_255
timestamp 1679581782
transform 1 0 25056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_262
timestamp 1679577901
transform 1 0 25728 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_266
timestamp 1677579658
transform 1 0 26112 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_271
timestamp 1677580104
transform 1 0 26592 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_277
timestamp 1677580104
transform 1 0 27168 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_293
timestamp 1677579658
transform 1 0 28704 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_298
timestamp 1677579658
transform 1 0 29184 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 30144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_315
timestamp 1679577901
transform 1 0 30816 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_319
timestamp 1677580104
transform 1 0 31200 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_325
timestamp 1677580104
transform 1 0 31776 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_331
timestamp 1679577901
transform 1 0 32352 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 33504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_364
timestamp 1677580104
transform 1 0 35520 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_379
timestamp 1679581782
transform 1 0 36960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_386
timestamp 1679581782
transform 1 0 37632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_393
timestamp 1679581782
transform 1 0 38304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_409
timestamp 1679581782
transform 1 0 39840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_416
timestamp 1679577901
transform 1 0 40512 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_420
timestamp 1677579658
transform 1 0 40896 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_425
timestamp 1679581782
transform 1 0 41376 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_432
timestamp 1677580104
transform 1 0 42048 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_471
timestamp 1677579658
transform 1 0 45792 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_499
timestamp 1677580104
transform 1 0 48480 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_501
timestamp 1677579658
transform 1 0 48672 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_507
timestamp 1677580104
transform 1 0 49248 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_539
timestamp 1677580104
transform 1 0 52320 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_25
timestamp 1677580104
transform 1 0 2976 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_31
timestamp 1679581782
transform 1 0 3552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_38
timestamp 1679581782
transform 1 0 4224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_45
timestamp 1679581782
transform 1 0 4896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_52
timestamp 1679581782
transform 1 0 5568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_59
timestamp 1679581782
transform 1 0 6240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_66
timestamp 1679581782
transform 1 0 6912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_73
timestamp 1679581782
transform 1 0 7584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_80
timestamp 1679581782
transform 1 0 8256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_87
timestamp 1679581782
transform 1 0 8928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_94
timestamp 1679581782
transform 1 0 9600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_101
timestamp 1679581782
transform 1 0 10272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_108
timestamp 1679581782
transform 1 0 10944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_115
timestamp 1679581782
transform 1 0 11616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_122
timestamp 1679581782
transform 1 0 12288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_129
timestamp 1679581782
transform 1 0 12960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_136
timestamp 1679581782
transform 1 0 13632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_143
timestamp 1679581782
transform 1 0 14304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_150
timestamp 1679581782
transform 1 0 14976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_157
timestamp 1679581782
transform 1 0 15648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_164
timestamp 1679581782
transform 1 0 16320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_171
timestamp 1679581782
transform 1 0 16992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_178
timestamp 1679581782
transform 1 0 17664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_185
timestamp 1679581782
transform 1 0 18336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_192
timestamp 1679581782
transform 1 0 19008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_199
timestamp 1679581782
transform 1 0 19680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_206
timestamp 1679581782
transform 1 0 20352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_213
timestamp 1679581782
transform 1 0 21024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_220
timestamp 1679581782
transform 1 0 21696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_227
timestamp 1679581782
transform 1 0 22368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_234
timestamp 1679581782
transform 1 0 23040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_241
timestamp 1679581782
transform 1 0 23712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_248
timestamp 1679581782
transform 1 0 24384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_255
timestamp 1679581782
transform 1 0 25056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_262
timestamp 1679581782
transform 1 0 25728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_269
timestamp 1679581782
transform 1 0 26400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_276
timestamp 1679581782
transform 1 0 27072 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_283
timestamp 1677580104
transform 1 0 27744 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_289
timestamp 1679581782
transform 1 0 28320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_296
timestamp 1679581782
transform 1 0 28992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_303
timestamp 1679577901
transform 1 0 29664 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_307
timestamp 1677580104
transform 1 0 30048 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_324
timestamp 1677579658
transform 1 0 31680 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_330
timestamp 1677580104
transform 1 0 32256 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_359
timestamp 1677580104
transform 1 0 35040 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_361
timestamp 1677579658
transform 1 0 35232 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_393
timestamp 1677580104
transform 1 0 38304 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_395
timestamp 1677579658
transform 1 0 38496 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_405
timestamp 1679581782
transform 1 0 39456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_448
timestamp 1679581782
transform 1 0 43584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_455
timestamp 1679581782
transform 1 0 44256 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_462
timestamp 1677579658
transform 1 0 44928 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_472
timestamp 1679577901
transform 1 0 45888 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_476
timestamp 1677579658
transform 1 0 46272 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_481
timestamp 1679581782
transform 1 0 46752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_488
timestamp 1679581782
transform 1 0 47424 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_513
timestamp 1677580104
transform 1 0 49824 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_515
timestamp 1677579658
transform 1 0 50016 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_533
timestamp 1677580104
transform 1 0 51744 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_4
timestamp 1679577901
transform 1 0 960 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_17
timestamp 1679581782
transform 1 0 2208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_24
timestamp 1679581782
transform 1 0 2880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_31
timestamp 1679581782
transform 1 0 3552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_38
timestamp 1679581782
transform 1 0 4224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_45
timestamp 1679581782
transform 1 0 4896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_52
timestamp 1679581782
transform 1 0 5568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_59
timestamp 1679581782
transform 1 0 6240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_66
timestamp 1679581782
transform 1 0 6912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_73
timestamp 1679581782
transform 1 0 7584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_80
timestamp 1679581782
transform 1 0 8256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_87
timestamp 1679581782
transform 1 0 8928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_94
timestamp 1679581782
transform 1 0 9600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_101
timestamp 1679581782
transform 1 0 10272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_108
timestamp 1679581782
transform 1 0 10944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_115
timestamp 1679581782
transform 1 0 11616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_122
timestamp 1679581782
transform 1 0 12288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_129
timestamp 1679581782
transform 1 0 12960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_136
timestamp 1679581782
transform 1 0 13632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_143
timestamp 1679581782
transform 1 0 14304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_150
timestamp 1679581782
transform 1 0 14976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_157
timestamp 1679581782
transform 1 0 15648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_164
timestamp 1679581782
transform 1 0 16320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_171
timestamp 1679581782
transform 1 0 16992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_178
timestamp 1679581782
transform 1 0 17664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_185
timestamp 1679581782
transform 1 0 18336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_192
timestamp 1679581782
transform 1 0 19008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_199
timestamp 1679581782
transform 1 0 19680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_206
timestamp 1679581782
transform 1 0 20352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_213
timestamp 1679581782
transform 1 0 21024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_220
timestamp 1679581782
transform 1 0 21696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_227
timestamp 1679581782
transform 1 0 22368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_234
timestamp 1679581782
transform 1 0 23040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_241
timestamp 1679581782
transform 1 0 23712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_248
timestamp 1679581782
transform 1 0 24384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_255
timestamp 1679581782
transform 1 0 25056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_262
timestamp 1679581782
transform 1 0 25728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_269
timestamp 1679581782
transform 1 0 26400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_276
timestamp 1679581782
transform 1 0 27072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_283
timestamp 1679577901
transform 1 0 27744 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_29_314
timestamp 1679577901
transform 1 0 30720 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_323
timestamp 1679581782
transform 1 0 31584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_347
timestamp 1679581782
transform 1 0 33888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_354
timestamp 1679581782
transform 1 0 34560 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_384
timestamp 1677580104
transform 1 0 37440 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_386
timestamp 1677579658
transform 1 0 37632 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_392
timestamp 1677580104
transform 1 0 38208 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_443
timestamp 1679581782
transform 1 0 43104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_450
timestamp 1679581782
transform 1 0 43776 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_457
timestamp 1677579658
transform 1 0 44448 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_463
timestamp 1679577901
transform 1 0 45024 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_476
timestamp 1677579658
transform 1 0 46272 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_504
timestamp 1677580104
transform 1 0 48960 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_506
timestamp 1677579658
transform 1 0 49152 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_534
timestamp 1679581782
transform 1 0 51840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_4
timestamp 1679577901
transform 1 0 960 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_8
timestamp 1677580104
transform 1 0 1344 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_18
timestamp 1679581782
transform 1 0 2304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_25
timestamp 1679581782
transform 1 0 2976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_32
timestamp 1679581782
transform 1 0 3648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_39
timestamp 1679581782
transform 1 0 4320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_46
timestamp 1679581782
transform 1 0 4992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_53
timestamp 1679581782
transform 1 0 5664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_60
timestamp 1679581782
transform 1 0 6336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_67
timestamp 1679581782
transform 1 0 7008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_74
timestamp 1679581782
transform 1 0 7680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_81
timestamp 1679581782
transform 1 0 8352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_88
timestamp 1679581782
transform 1 0 9024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_95
timestamp 1679581782
transform 1 0 9696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_102
timestamp 1679581782
transform 1 0 10368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_109
timestamp 1679581782
transform 1 0 11040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_116
timestamp 1679581782
transform 1 0 11712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_123
timestamp 1679581782
transform 1 0 12384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_130
timestamp 1679581782
transform 1 0 13056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_137
timestamp 1679581782
transform 1 0 13728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_144
timestamp 1679581782
transform 1 0 14400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_151
timestamp 1679581782
transform 1 0 15072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_158
timestamp 1679581782
transform 1 0 15744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_165
timestamp 1679581782
transform 1 0 16416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_172
timestamp 1679581782
transform 1 0 17088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_179
timestamp 1679581782
transform 1 0 17760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_186
timestamp 1679581782
transform 1 0 18432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_193
timestamp 1679581782
transform 1 0 19104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_200
timestamp 1679581782
transform 1 0 19776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_207
timestamp 1679581782
transform 1 0 20448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_214
timestamp 1679581782
transform 1 0 21120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_221
timestamp 1679581782
transform 1 0 21792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_228
timestamp 1679581782
transform 1 0 22464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_235
timestamp 1679581782
transform 1 0 23136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_242
timestamp 1679581782
transform 1 0 23808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_249
timestamp 1679581782
transform 1 0 24480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_256
timestamp 1679581782
transform 1 0 25152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_263
timestamp 1679581782
transform 1 0 25824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_270
timestamp 1679581782
transform 1 0 26496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_277
timestamp 1679581782
transform 1 0 27168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_284
timestamp 1679581782
transform 1 0 27840 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_291
timestamp 1677579658
transform 1 0 28512 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_296
timestamp 1679581782
transform 1 0 28992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_303
timestamp 1679581782
transform 1 0 29664 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_310
timestamp 1677580104
transform 1 0 30336 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_312
timestamp 1677579658
transform 1 0 30528 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_318
timestamp 1677580104
transform 1 0 31104 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_320
timestamp 1677579658
transform 1 0 31296 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_325
timestamp 1677579658
transform 1 0 31776 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_336
timestamp 1677580104
transform 1 0 32832 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_365
timestamp 1677580104
transform 1 0 35616 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_385
timestamp 1679581782
transform 1 0 37536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_392
timestamp 1679577901
transform 1 0 38208 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_396
timestamp 1677580104
transform 1 0 38592 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_408
timestamp 1679581782
transform 1 0 39744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_446
timestamp 1679577901
transform 1 0 43392 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_450
timestamp 1677579658
transform 1 0 43776 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_461
timestamp 1677579658
transform 1 0 44832 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_476
timestamp 1679577901
transform 1 0 46272 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_480
timestamp 1677580104
transform 1 0 46656 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_486
timestamp 1679581782
transform 1 0 47232 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_530
timestamp 1677580104
transform 1 0 51456 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_559
timestamp 1679577901
transform 1 0 54240 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_563
timestamp 1677579658
transform 1 0 54624 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_584
timestamp 1677579658
transform 1 0 56640 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_588
timestamp 1677580104
transform 1 0 57024 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_593
timestamp 1677579658
transform 1 0 57504 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_597
timestamp 1677579658
transform 1 0 57888 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_601
timestamp 1677579658
transform 1 0 58272 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_605
timestamp 1677580104
transform 1 0 58656 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_610
timestamp 1677579658
transform 1 0 59136 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_614
timestamp 1677579658
transform 1 0 59520 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_618
timestamp 1677579658
transform 1 0 59904 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_622
timestamp 1677579658
transform 1 0 60288 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_626
timestamp 1677579658
transform 1 0 60672 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_630
timestamp 1677580104
transform 1 0 61056 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_635
timestamp 1677579658
transform 1 0 61536 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_639
timestamp 1677579658
transform 1 0 61920 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_643
timestamp 1677579658
transform 1 0 62304 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_647
timestamp 1677579658
transform 1 0 62688 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_651
timestamp 1677579658
transform 1 0 63072 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_655
timestamp 1677580104
transform 1 0 63456 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_660
timestamp 1677579658
transform 1 0 63936 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_664
timestamp 1677579658
transform 1 0 64320 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_668
timestamp 1677579658
transform 1 0 64704 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_672
timestamp 1677579658
transform 1 0 65088 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_676
timestamp 1677580104
transform 1 0 65472 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_681
timestamp 1677579658
transform 1 0 65952 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_685
timestamp 1677579658
transform 1 0 66336 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_689
timestamp 1677579658
transform 1 0 66720 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_693
timestamp 1677579658
transform 1 0 67104 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_697
timestamp 1677580104
transform 1 0 67488 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_702
timestamp 1677579658
transform 1 0 67968 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_706
timestamp 1677579658
transform 1 0 68352 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_710
timestamp 1677579658
transform 1 0 68736 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_714
timestamp 1677579658
transform 1 0 69120 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_718
timestamp 1677580104
transform 1 0 69504 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_723
timestamp 1677579658
transform 1 0 69984 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_727
timestamp 1677579658
transform 1 0 70368 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_731
timestamp 1677579658
transform 1 0 70752 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_735
timestamp 1677579658
transform 1 0 71136 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_739
timestamp 1677579658
transform 1 0 71520 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_743
timestamp 1677579658
transform 1 0 71904 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_747
timestamp 1677579658
transform 1 0 72288 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_751
timestamp 1677579658
transform 1 0 72672 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_755
timestamp 1677580104
transform 1 0 73056 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_760
timestamp 1677579658
transform 1 0 73536 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_764
timestamp 1677579658
transform 1 0 73920 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_768
timestamp 1677579658
transform 1 0 74304 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_772
timestamp 1677579658
transform 1 0 74688 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_776
timestamp 1677579658
transform 1 0 75072 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_780
timestamp 1677579658
transform 1 0 75456 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_784
timestamp 1677580104
transform 1 0 75840 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_789
timestamp 1679577901
transform 1 0 76320 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_793
timestamp 1677579658
transform 1 0 76704 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_806
timestamp 1677579658
transform 1 0 77952 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_810
timestamp 1677579658
transform 1 0 78336 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_11
timestamp 1679581782
transform 1 0 1632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_25
timestamp 1679581782
transform 1 0 2976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_32
timestamp 1679581782
transform 1 0 3648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_39
timestamp 1679581782
transform 1 0 4320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_46
timestamp 1679581782
transform 1 0 4992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_53
timestamp 1679581782
transform 1 0 5664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_60
timestamp 1679581782
transform 1 0 6336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_67
timestamp 1679581782
transform 1 0 7008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_74
timestamp 1679581782
transform 1 0 7680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_81
timestamp 1679581782
transform 1 0 8352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_88
timestamp 1679581782
transform 1 0 9024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_95
timestamp 1679581782
transform 1 0 9696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_102
timestamp 1679581782
transform 1 0 10368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_109
timestamp 1679581782
transform 1 0 11040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_116
timestamp 1679581782
transform 1 0 11712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_123
timestamp 1679581782
transform 1 0 12384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_130
timestamp 1679581782
transform 1 0 13056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_137
timestamp 1679581782
transform 1 0 13728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_144
timestamp 1679581782
transform 1 0 14400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_151
timestamp 1679581782
transform 1 0 15072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_158
timestamp 1679581782
transform 1 0 15744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_165
timestamp 1679581782
transform 1 0 16416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_172
timestamp 1679581782
transform 1 0 17088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_179
timestamp 1679581782
transform 1 0 17760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_186
timestamp 1679581782
transform 1 0 18432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_193
timestamp 1679581782
transform 1 0 19104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_200
timestamp 1679581782
transform 1 0 19776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_207
timestamp 1679581782
transform 1 0 20448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_214
timestamp 1679581782
transform 1 0 21120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_221
timestamp 1679581782
transform 1 0 21792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_228
timestamp 1679581782
transform 1 0 22464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_235
timestamp 1679581782
transform 1 0 23136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_242
timestamp 1679581782
transform 1 0 23808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_249
timestamp 1679581782
transform 1 0 24480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_256
timestamp 1679581782
transform 1 0 25152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_263
timestamp 1679581782
transform 1 0 25824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_270
timestamp 1679581782
transform 1 0 26496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_277
timestamp 1679581782
transform 1 0 27168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_284
timestamp 1679581782
transform 1 0 27840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_291
timestamp 1679581782
transform 1 0 28512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_298
timestamp 1679577901
transform 1 0 29184 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_302
timestamp 1677580104
transform 1 0 29568 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_336
timestamp 1679581782
transform 1 0 32832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_343
timestamp 1679581782
transform 1 0 33504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679581782
transform 1 0 34176 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_357
timestamp 1677580104
transform 1 0 34848 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_386
timestamp 1679581782
transform 1 0 37632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_393
timestamp 1679581782
transform 1 0 38304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_423
timestamp 1679581782
transform 1 0 41184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_430
timestamp 1679577901
transform 1 0 41856 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_466
timestamp 1679581782
transform 1 0 45312 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_473
timestamp 1677579658
transform 1 0 45984 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_493
timestamp 1679577901
transform 1 0 47904 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_497
timestamp 1677579658
transform 1 0 48288 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_502
timestamp 1679581782
transform 1 0 48768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_509
timestamp 1679577901
transform 1 0 49440 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_513
timestamp 1677579658
transform 1 0 49824 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_523
timestamp 1677580104
transform 1 0 50784 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_525
timestamp 1677579658
transform 1 0 50976 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_530
timestamp 1679577901
transform 1 0 51456 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_534
timestamp 1677580104
transform 1 0 51840 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_545
timestamp 1679581782
transform 1 0 52896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_552
timestamp 1679581782
transform 1 0 53568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_559
timestamp 1679581782
transform 1 0 54240 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_566
timestamp 1677579658
transform 1 0 54912 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_594
timestamp 1679577901
transform 1 0 57600 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_603
timestamp 1677580104
transform 1 0 58464 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_631
timestamp 1679581782
transform 1 0 61152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_638
timestamp 1679581782
transform 1 0 61824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_645
timestamp 1679581782
transform 1 0 62496 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_652
timestamp 1677580104
transform 1 0 63168 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_654
timestamp 1677579658
transform 1 0 63360 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_672
timestamp 1679581782
transform 1 0 65088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_679
timestamp 1679581782
transform 1 0 65760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_686
timestamp 1679581782
transform 1 0 66432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_693
timestamp 1679577901
transform 1 0 67104 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_697
timestamp 1677579658
transform 1 0 67488 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_711
timestamp 1679581782
transform 1 0 68832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_718
timestamp 1679581782
transform 1 0 69504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_725
timestamp 1679577901
transform 1 0 70176 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_729
timestamp 1677579658
transform 1 0 70560 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_743
timestamp 1679581782
transform 1 0 71904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_750
timestamp 1679581782
transform 1 0 72576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_757
timestamp 1679581782
transform 1 0 73248 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_764
timestamp 1677580104
transform 1 0 73920 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_766
timestamp 1677579658
transform 1 0 74112 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_772
timestamp 1679577901
transform 1 0 74688 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_776
timestamp 1677580104
transform 1 0 75072 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_788
timestamp 1677580104
transform 1 0 76224 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_794
timestamp 1677580104
transform 1 0 76800 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_796
timestamp 1677579658
transform 1 0 76992 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_801
timestamp 1679581782
transform 1 0 77472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_808
timestamp 1679581782
transform 1 0 78144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_815
timestamp 1679581782
transform 1 0 78816 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_822
timestamp 1677579658
transform 1 0 79488 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1679581782
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_39
timestamp 1679581782
transform 1 0 4320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 4992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 5664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_60
timestamp 1679581782
transform 1 0 6336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679581782
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679581782
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679581782
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679581782
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_109
timestamp 1679581782
transform 1 0 11040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_116
timestamp 1679581782
transform 1 0 11712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_123
timestamp 1679581782
transform 1 0 12384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_130
timestamp 1679581782
transform 1 0 13056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_137
timestamp 1679581782
transform 1 0 13728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_144
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_158
timestamp 1679581782
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679581782
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679581782
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679581782
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679581782
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679581782
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679581782
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679581782
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_221
timestamp 1679581782
transform 1 0 21792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679581782
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679581782
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_249
timestamp 1679581782
transform 1 0 24480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_256
timestamp 1679581782
transform 1 0 25152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_263
timestamp 1679581782
transform 1 0 25824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_270
timestamp 1679581782
transform 1 0 26496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_277
timestamp 1679581782
transform 1 0 27168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_284
timestamp 1679581782
transform 1 0 27840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_291
timestamp 1679581782
transform 1 0 28512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_298
timestamp 1679581782
transform 1 0 29184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_305
timestamp 1679577901
transform 1 0 29856 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_313
timestamp 1679581782
transform 1 0 30624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_320
timestamp 1679577901
transform 1 0 31296 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_324
timestamp 1677580104
transform 1 0 31680 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_331
timestamp 1677579658
transform 1 0 32352 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_336
timestamp 1677580104
transform 1 0 32832 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_338
timestamp 1677579658
transform 1 0 33024 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_344
timestamp 1679577901
transform 1 0 33600 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_348
timestamp 1677580104
transform 1 0 33984 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_360
timestamp 1677579658
transform 1 0 35136 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_370
timestamp 1677580104
transform 1 0 36096 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_375
timestamp 1679577901
transform 1 0 36576 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_379
timestamp 1677580104
transform 1 0 36960 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_421
timestamp 1677580104
transform 1 0 40992 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_423
timestamp 1677579658
transform 1 0 41184 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_428
timestamp 1679581782
transform 1 0 41664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_435
timestamp 1679577901
transform 1 0 42336 0 1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_32_443
timestamp 1679577901
transform 1 0 43104 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_447
timestamp 1677579658
transform 1 0 43488 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_479
timestamp 1677579658
transform 1 0 46560 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_511
timestamp 1679581782
transform 1 0 49632 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_518
timestamp 1677580104
transform 1 0 50304 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_566
timestamp 1679577901
transform 1 0 54912 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_578
timestamp 1679581782
transform 1 0 56064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_585
timestamp 1679581782
transform 1 0 56736 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_619
timestamp 1677579658
transform 1 0 60000 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_647
timestamp 1677580104
transform 1 0 62688 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_649
timestamp 1677579658
transform 1 0 62880 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_687
timestamp 1679577901
transform 1 0 66528 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_728
timestamp 1677579658
transform 1 0 70464 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_819
timestamp 1679577901
transform 1 0 79200 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_4
timestamp 1679581782
transform 1 0 960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_11
timestamp 1679581782
transform 1 0 1632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_18
timestamp 1679581782
transform 1 0 2304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_25
timestamp 1679581782
transform 1 0 2976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_32
timestamp 1679581782
transform 1 0 3648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_39
timestamp 1679581782
transform 1 0 4320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679581782
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_53
timestamp 1679581782
transform 1 0 5664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_60
timestamp 1679581782
transform 1 0 6336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_67
timestamp 1679581782
transform 1 0 7008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_74
timestamp 1679581782
transform 1 0 7680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_81
timestamp 1679581782
transform 1 0 8352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_88
timestamp 1679581782
transform 1 0 9024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_95
timestamp 1679581782
transform 1 0 9696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_102
timestamp 1679581782
transform 1 0 10368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_109
timestamp 1679581782
transform 1 0 11040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_116
timestamp 1679581782
transform 1 0 11712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_123
timestamp 1679581782
transform 1 0 12384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_130
timestamp 1679581782
transform 1 0 13056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_137
timestamp 1679581782
transform 1 0 13728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_144
timestamp 1679581782
transform 1 0 14400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_151
timestamp 1679581782
transform 1 0 15072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_158
timestamp 1679581782
transform 1 0 15744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_165
timestamp 1679581782
transform 1 0 16416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_172
timestamp 1679581782
transform 1 0 17088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_179
timestamp 1679581782
transform 1 0 17760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_186
timestamp 1679581782
transform 1 0 18432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_193
timestamp 1679581782
transform 1 0 19104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_200
timestamp 1679581782
transform 1 0 19776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_207
timestamp 1679581782
transform 1 0 20448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_214
timestamp 1679581782
transform 1 0 21120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_221
timestamp 1679581782
transform 1 0 21792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_228
timestamp 1679581782
transform 1 0 22464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_235
timestamp 1679581782
transform 1 0 23136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_242
timestamp 1679581782
transform 1 0 23808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_249
timestamp 1679581782
transform 1 0 24480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_256
timestamp 1679581782
transform 1 0 25152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_263
timestamp 1679581782
transform 1 0 25824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_270
timestamp 1679581782
transform 1 0 26496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_277
timestamp 1679581782
transform 1 0 27168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_284
timestamp 1679581782
transform 1 0 27840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_291
timestamp 1679581782
transform 1 0 28512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_298
timestamp 1679581782
transform 1 0 29184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_305
timestamp 1679581782
transform 1 0 29856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_312
timestamp 1679581782
transform 1 0 30528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_319
timestamp 1679581782
transform 1 0 31200 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_368
timestamp 1677580104
transform 1 0 35904 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_370
timestamp 1677579658
transform 1 0 36096 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_379
timestamp 1679581782
transform 1 0 36960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_390
timestamp 1679581782
transform 1 0 38016 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_397
timestamp 1677579658
transform 1 0 38688 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_412
timestamp 1677580104
transform 1 0 40128 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_422
timestamp 1677580104
transform 1 0 41088 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_429
timestamp 1679577901
transform 1 0 41760 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_437
timestamp 1679581782
transform 1 0 42528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_444
timestamp 1679577901
transform 1 0 43200 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_448
timestamp 1677580104
transform 1 0 43584 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_482
timestamp 1677580104
transform 1 0 46848 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_484
timestamp 1677579658
transform 1 0 47040 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_538
timestamp 1677580104
transform 1 0 52224 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_548
timestamp 1679581782
transform 1 0 53184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_555
timestamp 1679581782
transform 1 0 53856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_562
timestamp 1679577901
transform 1 0 54528 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_590
timestamp 1679581782
transform 1 0 57216 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_610
timestamp 1677579658
transform 1 0 59136 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_632
timestamp 1677580104
transform 1 0 61248 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_634
timestamp 1677579658
transform 1 0 61440 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_672
timestamp 1677580104
transform 1 0 65088 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_679
timestamp 1679577901
transform 1 0 65760 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_687
timestamp 1679577901
transform 1 0 66528 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_691
timestamp 1677580104
transform 1 0 66912 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_707
timestamp 1677579658
transform 1 0 68448 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_712
timestamp 1677580104
transform 1 0 68928 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_714
timestamp 1677579658
transform 1 0 69120 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_720
timestamp 1679581782
transform 1 0 69696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_745
timestamp 1679581782
transform 1 0 72096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_752
timestamp 1679577901
transform 1 0 72768 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_760
timestamp 1679577901
transform 1 0 73536 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_764
timestamp 1677580104
transform 1 0 73920 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_781
timestamp 1679581782
transform 1 0 75552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_788
timestamp 1679577901
transform 1 0 76224 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_792
timestamp 1677579658
transform 1 0 76608 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_798
timestamp 1679581782
transform 1 0 77184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_805
timestamp 1679581782
transform 1 0 77856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_812
timestamp 1679581782
transform 1 0 78528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_819
timestamp 1679577901
transform 1 0 79200 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679581782
transform 1 0 10656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679581782
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679581782
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679581782
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679581782
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679581782
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679581782
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679581782
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679581782
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679581782
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679581782
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679581782
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679581782
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679581782
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679581782
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679581782
transform 1 0 28800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679581782
transform 1 0 29472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679581782
transform 1 0 30144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679581782
transform 1 0 30816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679581782
transform 1 0 31488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679581782
transform 1 0 32160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679581782
transform 1 0 32832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679581782
transform 1 0 33504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679581782
transform 1 0 34176 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_357
timestamp 1677579658
transform 1 0 34848 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_362
timestamp 1677580104
transform 1 0 35328 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_364
timestamp 1677579658
transform 1 0 35520 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_396
timestamp 1679577901
transform 1 0 38592 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_400
timestamp 1677579658
transform 1 0 38976 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_455
timestamp 1679577901
transform 1 0 44256 0 1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_34_511
timestamp 1679577901
transform 1 0 49632 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_515
timestamp 1677579658
transform 1 0 50016 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679581782
transform 1 0 52320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679581782
transform 1 0 52992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_553
timestamp 1679577901
transform 1 0 53664 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_557
timestamp 1677579658
transform 1 0 54048 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_585
timestamp 1679581782
transform 1 0 56736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_592
timestamp 1679577901
transform 1 0 57408 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_596
timestamp 1677579658
transform 1 0 57792 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_605
timestamp 1677579658
transform 1 0 58656 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_611
timestamp 1677579658
transform 1 0 59232 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_634
timestamp 1679577901
transform 1 0 61440 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_638
timestamp 1677580104
transform 1 0 61824 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679581782
transform 1 0 62400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679581782
transform 1 0 63072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_663
timestamp 1679581782
transform 1 0 64224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_670
timestamp 1679581782
transform 1 0 64896 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_704
timestamp 1677579658
transform 1 0 68160 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_749
timestamp 1679577901
transform 1 0 72480 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_753
timestamp 1677579658
transform 1 0 72864 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_28
timestamp 1679577901
transform 1 0 3264 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_385
timestamp 1677580104
transform 1 0 37536 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_419
timestamp 1677580104
transform 1 0 40800 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_429
timestamp 1679581782
transform 1 0 41760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_436
timestamp 1679581782
transform 1 0 42432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_443
timestamp 1679577901
transform 1 0 43104 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_496
timestamp 1679577901
transform 1 0 48192 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_500
timestamp 1677580104
transform 1 0 48576 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_529
timestamp 1677579658
transform 1 0 51360 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_567
timestamp 1677579658
transform 1 0 55008 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_582
timestamp 1679581782
transform 1 0 56448 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_589
timestamp 1677579658
transform 1 0 57120 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_622
timestamp 1677580104
transform 1 0 60288 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_651
timestamp 1679577901
transform 1 0 63072 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_655
timestamp 1677580104
transform 1 0 63456 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_662
timestamp 1679577901
transform 1 0 64128 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_666
timestamp 1677580104
transform 1 0 64512 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_681
timestamp 1677580104
transform 1 0 65952 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_687
timestamp 1679581782
transform 1 0 66528 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_694
timestamp 1677579658
transform 1 0 67200 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_699
timestamp 1679581782
transform 1 0 67680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_706
timestamp 1679581782
transform 1 0 68352 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_713
timestamp 1677579658
transform 1 0 69024 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_728
timestamp 1677579658
transform 1 0 70464 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_746
timestamp 1679581782
transform 1 0 72192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_753
timestamp 1679577901
transform 1 0 72864 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_757
timestamp 1677580104
transform 1 0 73248 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_763
timestamp 1679581782
transform 1 0 73824 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_770
timestamp 1677580104
transform 1 0 74496 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_772
timestamp 1677579658
transform 1 0 74688 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_778
timestamp 1677579658
transform 1 0 75264 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_784
timestamp 1679581782
transform 1 0 75840 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_791
timestamp 1677579658
transform 1 0 76512 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_796
timestamp 1677579658
transform 1 0 76992 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_805
timestamp 1679581782
transform 1 0 77856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_812
timestamp 1679581782
transform 1 0 78528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_819
timestamp 1679577901
transform 1 0 79200 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_399
timestamp 1679577901
transform 1 0 38880 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_403
timestamp 1677580104
transform 1 0 39264 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_418
timestamp 1677580104
transform 1 0 40704 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_420
timestamp 1677579658
transform 1 0 40896 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_457
timestamp 1677579658
transform 1 0 44448 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_477
timestamp 1677580104
transform 1 0 46368 0 1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_483
timestamp 1679577901
transform 1 0 46944 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_487
timestamp 1677580104
transform 1 0 47328 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_493
timestamp 1679581782
transform 1 0 47904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_500
timestamp 1679581782
transform 1 0 48576 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_511
timestamp 1677580104
transform 1 0 49632 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_513
timestamp 1677579658
transform 1 0 49824 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_524
timestamp 1677580104
transform 1 0 50880 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_530
timestamp 1677579658
transform 1 0 51456 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_535
timestamp 1677579658
transform 1 0 51936 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679581782
transform 1 0 57024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_599
timestamp 1679577901
transform 1 0 58080 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_603
timestamp 1677580104
transform 1 0 58464 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_618
timestamp 1677580104
transform 1 0 59904 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_637
timestamp 1677579658
transform 1 0 61728 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_675
timestamp 1677580104
transform 1 0 65376 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_677
timestamp 1677579658
transform 1 0 65568 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_705
timestamp 1679581782
transform 1 0 68256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_712
timestamp 1679581782
transform 1 0 68928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_719
timestamp 1679577901
transform 1 0 69600 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_723
timestamp 1677579658
transform 1 0 69984 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_734
timestamp 1677580104
transform 1 0 71040 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_736
timestamp 1677579658
transform 1 0 71232 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_764
timestamp 1679581782
transform 1 0 73920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_771
timestamp 1679577901
transform 1 0 74592 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_775
timestamp 1677580104
transform 1 0 74976 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_782
timestamp 1679581782
transform 1 0 75648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_789
timestamp 1679577901
transform 1 0 76320 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_802
timestamp 1679581782
transform 1 0 77568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_809
timestamp 1679581782
transform 1 0 78240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_816
timestamp 1679581782
transform 1 0 78912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_392
timestamp 1677580104
transform 1 0 38208 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_440
timestamp 1679581782
transform 1 0 42816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_447
timestamp 1679581782
transform 1 0 43488 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_454
timestamp 1677580104
transform 1 0 44160 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_456
timestamp 1677579658
transform 1 0 44352 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_461
timestamp 1677580104
transform 1 0 44832 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_468
timestamp 1677579658
transform 1 0 45504 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_479
timestamp 1679581782
transform 1 0 46560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_486
timestamp 1679581782
transform 1 0 47232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_493
timestamp 1679581782
transform 1 0 47904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_500
timestamp 1679581782
transform 1 0 48576 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_507
timestamp 1677579658
transform 1 0 49248 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_521
timestamp 1677580104
transform 1 0 50592 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_528
timestamp 1679581782
transform 1 0 51264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_535
timestamp 1679581782
transform 1 0 51936 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_542
timestamp 1677580104
transform 1 0 52608 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_576
timestamp 1677580104
transform 1 0 55872 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_605
timestamp 1679577901
transform 1 0 58656 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_609
timestamp 1677579658
transform 1 0 59040 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_619
timestamp 1677580104
transform 1 0 60000 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_621
timestamp 1677579658
transform 1 0 60192 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_631
timestamp 1679581782
transform 1 0 61152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_638
timestamp 1679577901
transform 1 0 61824 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_642
timestamp 1677579658
transform 1 0 62208 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_647
timestamp 1679577901
transform 1 0 62688 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_651
timestamp 1677580104
transform 1 0 63072 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_663
timestamp 1679581782
transform 1 0 64224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_670
timestamp 1679581782
transform 1 0 64896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_682
timestamp 1679581782
transform 1 0 66048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_689
timestamp 1679577901
transform 1 0 66720 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_693
timestamp 1677579658
transform 1 0 67104 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_746
timestamp 1679581782
transform 1 0 72192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_753
timestamp 1679577901
transform 1 0 72864 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_757
timestamp 1677579658
transform 1 0 73248 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_795
timestamp 1677579658
transform 1 0 76896 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_403
timestamp 1679581782
transform 1 0 39264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_436
timestamp 1679581782
transform 1 0 42432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_443
timestamp 1679577901
transform 1 0 43104 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_505
timestamp 1677580104
transform 1 0 49056 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_526
timestamp 1677579658
transform 1 0 51072 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_554
timestamp 1679581782
transform 1 0 53760 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_561
timestamp 1677580104
transform 1 0 54432 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_563
timestamp 1677579658
transform 1 0 54624 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_569
timestamp 1679577901
transform 1 0 55200 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_577
timestamp 1677580104
transform 1 0 55968 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_587
timestamp 1679581782
transform 1 0 56928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_594
timestamp 1679577901
transform 1 0 57600 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_598
timestamp 1677580104
transform 1 0 57984 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_604
timestamp 1677580104
transform 1 0 58560 0 1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_38_662
timestamp 1679577901
transform 1 0 64128 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_666
timestamp 1677579658
transform 1 0 64512 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_708
timestamp 1679577901
transform 1 0 68544 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_712
timestamp 1677579658
transform 1 0 68928 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_736
timestamp 1677580104
transform 1 0 71232 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_747
timestamp 1679581782
transform 1 0 72288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_754
timestamp 1679581782
transform 1 0 72960 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_761
timestamp 1677580104
transform 1 0 73632 0 1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_38_767
timestamp 1679577901
transform 1 0 74208 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_771
timestamp 1677580104
transform 1 0 74592 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_787
timestamp 1677580104
transform 1 0 76128 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_789
timestamp 1677579658
transform 1 0 76320 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_794
timestamp 1677580104
transform 1 0 76800 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_805
timestamp 1679581782
transform 1 0 77856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_812
timestamp 1679581782
transform 1 0 78528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_819
timestamp 1679577901
transform 1 0 79200 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_413
timestamp 1677580104
transform 1 0 40224 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_415
timestamp 1677579658
transform 1 0 40416 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_424
timestamp 1679581782
transform 1 0 41280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_431
timestamp 1679577901
transform 1 0 41952 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_448
timestamp 1677580104
transform 1 0 43584 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_450
timestamp 1677579658
transform 1 0 43776 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_460
timestamp 1677579658
transform 1 0 44736 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_466
timestamp 1679577901
transform 1 0 45312 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_470
timestamp 1677579658
transform 1 0 45696 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_480
timestamp 1677580104
transform 1 0 46656 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_482
timestamp 1677579658
transform 1 0 46848 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_487
timestamp 1679581782
transform 1 0 47328 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_521
timestamp 1677579658
transform 1 0 50592 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_542
timestamp 1679577901
transform 1 0 52608 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_546
timestamp 1677580104
transform 1 0 52992 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_552
timestamp 1679581782
transform 1 0 53568 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_559
timestamp 1677580104
transform 1 0 54240 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_585
timestamp 1679581782
transform 1 0 56736 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_592
timestamp 1677580104
transform 1 0 57408 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_594
timestamp 1677579658
transform 1 0 57600 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_638
timestamp 1679581782
transform 1 0 61824 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_645
timestamp 1677579658
transform 1 0 62496 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_678
timestamp 1677580104
transform 1 0 65664 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_684
timestamp 1677580104
transform 1 0 66240 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_690
timestamp 1679581782
transform 1 0 66816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_697
timestamp 1679581782
transform 1 0 67488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_768
timestamp 1679577901
transform 1 0 74304 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_772
timestamp 1677579658
transform 1 0 74688 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_783
timestamp 1677580104
transform 1 0 75744 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_785
timestamp 1677579658
transform 1 0 75936 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_406
timestamp 1679577901
transform 1 0 39552 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_410
timestamp 1677579658
transform 1 0 39936 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_453
timestamp 1679581782
transform 1 0 44064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_460
timestamp 1679581782
transform 1 0 44736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_467
timestamp 1679581782
transform 1 0 45408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_474
timestamp 1679581782
transform 1 0 46080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_481
timestamp 1679581782
transform 1 0 46752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_488
timestamp 1679581782
transform 1 0 47424 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_504
timestamp 1677580104
transform 1 0 48960 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_535
timestamp 1679581782
transform 1 0 51936 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_542
timestamp 1677579658
transform 1 0 52608 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_570
timestamp 1677580104
transform 1 0 55296 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_576
timestamp 1677580104
transform 1 0 55872 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_605
timestamp 1679581782
transform 1 0 58656 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_612
timestamp 1677580104
transform 1 0 59328 0 1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_40_619
timestamp 1679577901
transform 1 0 60000 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_627
timestamp 1677580104
transform 1 0 60768 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_629
timestamp 1677579658
transform 1 0 60960 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_634
timestamp 1679581782
transform 1 0 61440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_641
timestamp 1679577901
transform 1 0 62112 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_655
timestamp 1677579658
transform 1 0 63456 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_660
timestamp 1679581782
transform 1 0 63936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_667
timestamp 1679581782
transform 1 0 64608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_674
timestamp 1679581782
transform 1 0 65280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_681
timestamp 1679577901
transform 1 0 65952 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_698
timestamp 1679581782
transform 1 0 67584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_705
timestamp 1679577901
transform 1 0 68256 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_709
timestamp 1677579658
transform 1 0 68640 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679581782
transform 1 0 69120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_721
timestamp 1679577901
transform 1 0 69792 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_725
timestamp 1677580104
transform 1 0 70176 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_736
timestamp 1677579658
transform 1 0 71232 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_741
timestamp 1679577901
transform 1 0 71712 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_745
timestamp 1677579658
transform 1 0 72096 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_750
timestamp 1679581782
transform 1 0 72576 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_757
timestamp 1677580104
transform 1 0 73248 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_759
timestamp 1677579658
transform 1 0 73440 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_787
timestamp 1679581782
transform 1 0 76128 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_794
timestamp 1677579658
transform 1 0 76800 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_799
timestamp 1677579658
transform 1 0 77280 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_808
timestamp 1679581782
transform 1 0 78144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_815
timestamp 1679581782
transform 1 0 78816 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_822
timestamp 1677579658
transform 1 0 79488 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_413
timestamp 1677580104
transform 1 0 40224 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_415
timestamp 1677579658
transform 1 0 40416 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_434
timestamp 1677579658
transform 1 0 42240 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_519
timestamp 1679581782
transform 1 0 50400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_553
timestamp 1679577901
transform 1 0 53664 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679581782
transform 1 0 55008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679581782
transform 1 0 55680 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_581
timestamp 1677580104
transform 1 0 56352 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_587
timestamp 1679581782
transform 1 0 56928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_594
timestamp 1679577901
transform 1 0 57600 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_598
timestamp 1677580104
transform 1 0 57984 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_619
timestamp 1677580104
transform 1 0 60000 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_621
timestamp 1677579658
transform 1 0 60192 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_667
timestamp 1679581782
transform 1 0 64608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_715
timestamp 1679577901
transform 1 0 69216 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_719
timestamp 1677579658
transform 1 0 69600 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_730
timestamp 1677579658
transform 1 0 70656 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_736
timestamp 1677580104
transform 1 0 71232 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_756
timestamp 1679581782
transform 1 0 73152 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_763
timestamp 1677580104
transform 1 0 73824 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_769
timestamp 1679581782
transform 1 0 74400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_776
timestamp 1679581782
transform 1 0 75072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_788
timestamp 1679577901
transform 1 0 76224 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_434
timestamp 1679577901
transform 1 0 42240 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_438
timestamp 1677579658
transform 1 0 42624 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_443
timestamp 1679581782
transform 1 0 43104 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_450
timestamp 1677579658
transform 1 0 43776 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679581782
transform 1 0 44256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679581782
transform 1 0 44928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_535
timestamp 1679581782
transform 1 0 51936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_542
timestamp 1679581782
transform 1 0 52608 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_549
timestamp 1677580104
transform 1 0 53280 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_551
timestamp 1677579658
transform 1 0 53472 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_557
timestamp 1679581782
transform 1 0 54048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_636
timestamp 1679581782
transform 1 0 61632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_648
timestamp 1679577901
transform 1 0 62784 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_679
timestamp 1677580104
transform 1 0 65760 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_691
timestamp 1679581782
transform 1 0 66912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_698
timestamp 1679581782
transform 1 0 67584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_705
timestamp 1679577901
transform 1 0 68256 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_709
timestamp 1677579658
transform 1 0 68640 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_742
timestamp 1677580104
transform 1 0 71808 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_744
timestamp 1677579658
transform 1 0 72000 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_813
timestamp 1679581782
transform 1 0 78624 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_820
timestamp 1677580104
transform 1 0 79296 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_822
timestamp 1677579658
transform 1 0 79488 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_469
timestamp 1679577901
transform 1 0 45600 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_482
timestamp 1679581782
transform 1 0 46848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_489
timestamp 1679581782
transform 1 0 47520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_496
timestamp 1679581782
transform 1 0 48192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_508
timestamp 1679581782
transform 1 0 49344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_515
timestamp 1679581782
transform 1 0 50016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_522
timestamp 1679581782
transform 1 0 50688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_529
timestamp 1679581782
transform 1 0 51360 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_536
timestamp 1677579658
transform 1 0 52032 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_43_574
timestamp 1679577901
transform 1 0 55680 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_582
timestamp 1679581782
transform 1 0 56448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_589
timestamp 1679581782
transform 1 0 57120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_596
timestamp 1679577901
transform 1 0 57792 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_600
timestamp 1677579658
transform 1 0 58176 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_614
timestamp 1679581782
transform 1 0 59520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_621
timestamp 1679581782
transform 1 0 60192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_628
timestamp 1679581782
transform 1 0 60864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_635
timestamp 1679577901
transform 1 0 61536 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_639
timestamp 1677580104
transform 1 0 61920 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_654
timestamp 1677580104
transform 1 0 63360 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_656
timestamp 1677579658
transform 1 0 63552 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_661
timestamp 1679581782
transform 1 0 64032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_668
timestamp 1679581782
transform 1 0 64704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_675
timestamp 1679581782
transform 1 0 65376 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_682
timestamp 1677579658
transform 1 0 66048 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_710
timestamp 1679581782
transform 1 0 68736 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_717
timestamp 1677580104
transform 1 0 69408 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_719
timestamp 1677579658
transform 1 0 69600 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_724
timestamp 1679581782
transform 1 0 70080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_731
timestamp 1679581782
transform 1 0 70752 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_738
timestamp 1677579658
transform 1 0 71424 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_752
timestamp 1679581782
transform 1 0 72768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_759
timestamp 1679581782
transform 1 0 73440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_766
timestamp 1679581782
transform 1 0 74112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_777
timestamp 1679577901
transform 1 0 75168 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_781
timestamp 1677579658
transform 1 0 75552 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_797
timestamp 1677579658
transform 1 0 77088 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_803
timestamp 1677579658
transform 1 0 77664 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_808
timestamp 1679581782
transform 1 0 78144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_815
timestamp 1679581782
transform 1 0 78816 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_822
timestamp 1677579658
transform 1 0 79488 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_469
timestamp 1677579658
transform 1 0 45600 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_501
timestamp 1679577901
transform 1 0 48672 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_505
timestamp 1677579658
transform 1 0 49056 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_518
timestamp 1677579658
transform 1 0 50304 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_529
timestamp 1677580104
transform 1 0 51360 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_535
timestamp 1677580104
transform 1 0 51936 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679581782
transform 1 0 52992 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_553
timestamp 1677580104
transform 1 0 53664 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_560
timestamp 1679577901
transform 1 0 54336 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_564
timestamp 1677580104
transform 1 0 54720 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_570
timestamp 1677580104
transform 1 0 55296 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_586
timestamp 1679577901
transform 1 0 56832 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_590
timestamp 1677580104
transform 1 0 57216 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_624
timestamp 1679581782
transform 1 0 60480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_631
timestamp 1679581782
transform 1 0 61152 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_643
timestamp 1677580104
transform 1 0 62304 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_677
timestamp 1679577901
transform 1 0 65568 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_681
timestamp 1677579658
transform 1 0 65952 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_700
timestamp 1677579658
transform 1 0 67776 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_705
timestamp 1679577901
transform 1 0 68256 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_709
timestamp 1677580104
transform 1 0 68640 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_738
timestamp 1677580104
transform 1 0 71424 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_772
timestamp 1679581782
transform 1 0 74688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_779
timestamp 1679577901
transform 1 0 75360 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_783
timestamp 1677580104
transform 1 0 75744 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_809
timestamp 1679581782
transform 1 0 78240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_816
timestamp 1679581782
transform 1 0 78912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_476
timestamp 1677580104
transform 1 0 46272 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_497
timestamp 1677579658
transform 1 0 48288 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_544
timestamp 1679581782
transform 1 0 52800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_551
timestamp 1679581782
transform 1 0 53472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_558
timestamp 1679577901
transform 1 0 54144 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_562
timestamp 1677579658
transform 1 0 54528 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_608
timestamp 1679581782
transform 1 0 58944 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_615
timestamp 1677579658
transform 1 0 59616 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_653
timestamp 1677580104
transform 1 0 63264 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_659
timestamp 1679581782
transform 1 0 63840 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_666
timestamp 1677579658
transform 1 0 64512 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_671
timestamp 1679581782
transform 1 0 64992 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_678
timestamp 1677579658
transform 1 0 65664 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_694
timestamp 1677580104
transform 1 0 67200 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_723
timestamp 1679577901
transform 1 0 69984 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_755
timestamp 1679581782
transform 1 0 73056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_762
timestamp 1679577901
transform 1 0 73728 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_793
timestamp 1677580104
transform 1 0 76704 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_795
timestamp 1677579658
transform 1 0 76896 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_497
timestamp 1679577901
transform 1 0 48288 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_501
timestamp 1677580104
transform 1 0 48672 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_507
timestamp 1679581782
transform 1 0 49248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_514
timestamp 1679581782
transform 1 0 49920 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_521
timestamp 1677579658
transform 1 0 50592 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_526
timestamp 1677579658
transform 1 0 51072 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_531
timestamp 1679577901
transform 1 0 51552 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_562
timestamp 1679581782
transform 1 0 54528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_569
timestamp 1679577901
transform 1 0 55200 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_573
timestamp 1677579658
transform 1 0 55584 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_587
timestamp 1679581782
transform 1 0 56928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_594
timestamp 1679581782
transform 1 0 57600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_601
timestamp 1679577901
transform 1 0 58272 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_605
timestamp 1677579658
transform 1 0 58656 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_610
timestamp 1679581782
transform 1 0 59136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_617
timestamp 1679577901
transform 1 0 59808 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_625
timestamp 1679581782
transform 1 0 60576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_642
timestamp 1679581782
transform 1 0 62208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_649
timestamp 1679581782
transform 1 0 62880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_656
timestamp 1679577901
transform 1 0 63552 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_660
timestamp 1677580104
transform 1 0 63936 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_698
timestamp 1679581782
transform 1 0 67584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_705
timestamp 1679581782
transform 1 0 68256 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_712
timestamp 1677580104
transform 1 0 68928 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_714
timestamp 1677579658
transform 1 0 69120 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_724
timestamp 1679581782
transform 1 0 70080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_731
timestamp 1679581782
transform 1 0 70752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_738
timestamp 1679577901
transform 1 0 71424 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_747
timestamp 1677580104
transform 1 0 72288 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_749
timestamp 1677579658
transform 1 0 72480 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_768
timestamp 1677580104
transform 1 0 74304 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_770
timestamp 1677579658
transform 1 0 74496 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_775
timestamp 1679581782
transform 1 0 74976 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_782
timestamp 1677580104
transform 1 0 75648 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_784
timestamp 1677579658
transform 1 0 75840 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_795
timestamp 1677579658
transform 1 0 76896 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_808
timestamp 1679581782
transform 1 0 78144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_815
timestamp 1679581782
transform 1 0 78816 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_822
timestamp 1677579658
transform 1 0 79488 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_592
timestamp 1679581782
transform 1 0 57408 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_618
timestamp 1677580104
transform 1 0 59904 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_625
timestamp 1679581782
transform 1 0 60576 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_632
timestamp 1677579658
transform 1 0 61248 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_643
timestamp 1679581782
transform 1 0 62304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_664
timestamp 1679581782
transform 1 0 64320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_671
timestamp 1679581782
transform 1 0 64992 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_705
timestamp 1677579658
transform 1 0 68256 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_723
timestamp 1679581782
transform 1 0 69984 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_730
timestamp 1677580104
transform 1 0 70656 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_560
timestamp 1679577901
transform 1 0 54336 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_564
timestamp 1677579658
transform 1 0 54720 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_569
timestamp 1677580104
transform 1 0 55200 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_608
timestamp 1677579658
transform 1 0 58944 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_690
timestamp 1677580104
transform 1 0 66816 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_711
timestamp 1677580104
transform 1 0 68832 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_740
timestamp 1679581782
transform 1 0 71616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_747
timestamp 1679577901
transform 1 0 72288 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_766
timestamp 1677579658
transform 1 0 74112 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_772
timestamp 1677580104
transform 1 0 74688 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_774
timestamp 1677579658
transform 1 0 74880 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_815
timestamp 1679581782
transform 1 0 78816 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_822
timestamp 1677579658
transform 1 0 79488 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_578
timestamp 1677580104
transform 1 0 56064 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_580
timestamp 1677579658
transform 1 0 56256 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_585
timestamp 1679577901
transform 1 0 56736 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_589
timestamp 1677579658
transform 1 0 57120 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_624
timestamp 1679581782
transform 1 0 60480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_631
timestamp 1679577901
transform 1 0 61152 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_635
timestamp 1677579658
transform 1 0 61536 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_640
timestamp 1679581782
transform 1 0 62016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_647
timestamp 1679581782
transform 1 0 62688 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_654
timestamp 1677579658
transform 1 0 63360 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_668
timestamp 1679581782
transform 1 0 64704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_675
timestamp 1679581782
transform 1 0 65376 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_682
timestamp 1677579658
transform 1 0 66048 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_687
timestamp 1679581782
transform 1 0 66528 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_694
timestamp 1677579658
transform 1 0 67200 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_707
timestamp 1677580104
transform 1 0 68448 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_714
timestamp 1677579658
transform 1 0 69120 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_745
timestamp 1679577901
transform 1 0 72096 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_749
timestamp 1677579658
transform 1 0 72480 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_763
timestamp 1677579658
transform 1 0 73824 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_768
timestamp 1679581782
transform 1 0 74304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_775
timestamp 1679581782
transform 1 0 74976 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_782
timestamp 1677580104
transform 1 0 75648 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_784
timestamp 1677579658
transform 1 0 75840 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_789
timestamp 1679577901
transform 1 0 76320 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_803
timestamp 1679581782
transform 1 0 77664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_810
timestamp 1679581782
transform 1 0 78336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_817
timestamp 1679577901
transform 1 0 79008 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_821
timestamp 1677580104
transform 1 0 79392 0 -1 38556
box -48 -56 240 834
use sg13g2_tiehi  heichips25_pudding_457
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_458
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_459
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_460
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_461
timestamp 1680000651
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_462
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_463
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 1344 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform -1 0 1344 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 1344 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
use analog_wires  wires
timestamp 0
transform 1 0 80000 0 1 800
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 16316 630 16756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 28316 630 28756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 40316 630 40756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 52316 630 52756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64316 630 64756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 76316 630 76756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 15076 712 15516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 27076 712 27516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 39076 712 39516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 51076 712 51516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63076 712 63516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 75076 712 75516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 99920 21586 100000 21726 0 FreeSans 640 0 0 0 i_in
port 4 nsew signal bidirectional
flabel metal3 s 99920 19949 100000 20089 0 FreeSans 640 0 0 0 i_out
port 5 nsew signal bidirectional
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 6 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 7 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 8 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 9 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 10 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 11 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 12 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 13 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 14 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 15 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 16 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 17 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 18 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 19 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 20 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 21 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 22 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 23 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 24 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 25 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 26 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 27 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 28 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 29 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 30 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 31 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 32 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 33 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 34 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 35 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 36 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 37 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 38 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 39 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 40 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 41 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 42 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 43 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 44 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 45 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 46 nsew signal output
rlabel via5 76620 22479 76620 22479 0 VGND
rlabel via5 75380 19603 75380 19603 0 VPWR
rlabel metal3 54048 17052 54048 17052 0 _0000_
rlabel metal2 64734 22764 64734 22764 0 _0001_
rlabel metal2 64342 22764 64342 22764 0 _0002_
rlabel metal2 63950 22764 63950 22764 0 _0003_
rlabel metal2 63565 22828 63565 22828 0 _0004_
rlabel metal2 63165 22828 63165 22828 0 _0005_
rlabel metal2 62765 22828 62765 22828 0 _0006_
rlabel metal2 62334 22764 62334 22764 0 _0007_
rlabel metal2 61942 22764 61942 22764 0 _0008_
rlabel metal2 61550 22764 61550 22764 0 _0009_
rlabel metal2 61165 22828 61165 22828 0 _0010_
rlabel metal2 58080 16758 58080 16758 0 _0011_
rlabel metal2 60765 22732 60765 22732 0 _0012_
rlabel metal2 60326 22764 60326 22764 0 _0013_
rlabel metal2 59934 22764 59934 22764 0 _0014_
rlabel metal2 59565 22828 59565 22828 0 _0015_
rlabel metal2 59165 22828 59165 22828 0 _0016_
rlabel metal2 58765 22828 58765 22828 0 _0017_
rlabel metal2 58270 22764 58270 22764 0 _0018_
rlabel metal2 57965 22828 57965 22828 0 _0019_
rlabel metal2 57565 22828 57565 22828 0 _0020_
rlabel metal2 57165 22828 57165 22828 0 _0021_
rlabel metal2 58368 16758 58368 16758 0 _0022_
rlabel metal2 56750 22764 56750 22764 0 _0023_
rlabel metal2 56365 22828 56365 22828 0 _0024_
rlabel metal2 55965 22828 55965 22828 0 _0025_
rlabel metal2 55565 22828 55565 22828 0 _0026_
rlabel metal2 55165 22828 55165 22828 0 _0027_
rlabel metal2 54765 22816 54765 22816 0 _0028_
rlabel metal2 54365 22828 54365 22828 0 _0029_
rlabel metal2 53965 22690 53965 22690 0 _0030_
rlabel metal2 58656 16758 58656 16758 0 _0031_
rlabel metal2 59136 16044 59136 16044 0 _0032_
rlabel metal2 59424 16086 59424 16086 0 _0033_
rlabel metal2 59904 16044 59904 16044 0 _0034_
rlabel metal2 60288 16464 60288 16464 0 _0035_
rlabel metal2 60672 16758 60672 16758 0 _0036_
rlabel metal2 61536 16758 61536 16758 0 _0037_
rlabel metal3 61968 16464 61968 16464 0 _0038_
rlabel metal2 54475 17763 54475 17763 0 _0039_
rlabel metal2 62400 16464 62400 16464 0 _0040_
rlabel metal2 62784 16002 62784 16002 0 _0041_
rlabel metal2 63072 16758 63072 16758 0 _0042_
rlabel metal2 63264 16758 63264 16758 0 _0043_
rlabel metal2 63648 16758 63648 16758 0 _0044_
rlabel metal2 63936 16758 63936 16758 0 _0045_
rlabel metal2 64320 16044 64320 16044 0 _0046_
rlabel metal2 64608 16800 64608 16800 0 _0047_
rlabel metal2 65088 16758 65088 16758 0 _0048_
rlabel metal2 65472 16758 65472 16758 0 _0049_
rlabel metal2 54528 16800 54528 16800 0 _0050_
rlabel metal2 65856 16758 65856 16758 0 _0051_
rlabel metal2 66336 16044 66336 16044 0 _0052_
rlabel metal2 66624 16800 66624 16800 0 _0053_
rlabel metal2 67104 16758 67104 16758 0 _0054_
rlabel metal2 67584 16464 67584 16464 0 _0055_
rlabel metal2 67872 16758 67872 16758 0 _0056_
rlabel metal2 68256 16758 68256 16758 0 _0057_
rlabel metal2 68736 16044 68736 16044 0 _0058_
rlabel metal2 69120 16758 69120 16758 0 _0059_
rlabel metal2 69504 16758 69504 16758 0 _0060_
rlabel metal2 54912 16758 54912 16758 0 _0061_
rlabel metal2 69888 16758 69888 16758 0 _0062_
rlabel metal2 70272 16758 70272 16758 0 _0063_
rlabel metal2 70656 16758 70656 16758 0 _0064_
rlabel metal2 71040 16758 71040 16758 0 _0065_
rlabel metal2 71424 16800 71424 16800 0 _0066_
rlabel metal2 71904 16758 71904 16758 0 _0067_
rlabel metal2 72288 16758 72288 16758 0 _0068_
rlabel metal2 72672 16758 72672 16758 0 _0069_
rlabel metal2 73056 16758 73056 16758 0 _0070_
rlabel metal2 73536 16758 73536 16758 0 _0071_
rlabel metal2 55488 16128 55488 16128 0 _0072_
rlabel metal2 73920 16044 73920 16044 0 _0073_
rlabel metal2 74304 16758 74304 16758 0 _0074_
rlabel metal2 74784 16464 74784 16464 0 _0075_
rlabel metal2 75072 16758 75072 16758 0 _0076_
rlabel metal2 75456 16758 75456 16758 0 _0077_
rlabel metal2 75840 16758 75840 16758 0 _0078_
rlabel metal2 76512 16758 76512 16758 0 _0079_
rlabel metal2 76896 16758 76896 16758 0 _0080_
rlabel metal2 77280 16758 77280 16758 0 _0081_
rlabel metal2 77568 16758 77568 16758 0 _0082_
rlabel metal2 55920 16464 55920 16464 0 _0083_
rlabel metal2 77952 16758 77952 16758 0 _0084_
rlabel metal2 78336 16758 78336 16758 0 _0085_
rlabel metal2 78720 16758 78720 16758 0 _0086_
rlabel metal2 79296 16800 79296 16800 0 _0087_
rlabel metal2 79165 22828 79165 22828 0 _0088_
rlabel metal2 78765 22828 78765 22828 0 _0089_
rlabel metal2 78350 22764 78350 22764 0 _0090_
rlabel metal2 77965 22828 77965 22828 0 _0091_
rlabel metal2 77565 22828 77565 22828 0 _0092_
rlabel metal2 77165 22828 77165 22828 0 _0093_
rlabel metal2 56256 16758 56256 16758 0 _0094_
rlabel metal2 76765 22828 76765 22828 0 _0095_
rlabel metal2 76342 22764 76342 22764 0 _0096_
rlabel metal2 75950 22764 75950 22764 0 _0097_
rlabel metal2 75565 22828 75565 22828 0 _0098_
rlabel metal2 75070 22764 75070 22764 0 _0099_
rlabel metal2 74765 22828 74765 22828 0 _0100_
rlabel metal2 74334 22764 74334 22764 0 _0101_
rlabel metal2 73942 22764 73942 22764 0 _0102_
rlabel metal2 73550 22764 73550 22764 0 _0103_
rlabel metal2 73165 22828 73165 22828 0 _0104_
rlabel metal2 56640 16590 56640 16590 0 _0105_
rlabel metal2 72670 22764 72670 22764 0 _0106_
rlabel metal2 72326 22764 72326 22764 0 _0107_
rlabel metal2 71934 22764 71934 22764 0 _0108_
rlabel metal2 71542 22764 71542 22764 0 _0109_
rlabel metal2 71150 22764 71150 22764 0 _0110_
rlabel metal2 70765 22828 70765 22828 0 _0111_
rlabel metal2 70365 22828 70365 22828 0 _0112_
rlabel metal2 69965 22828 69965 22828 0 _0113_
rlabel metal2 69534 22764 69534 22764 0 _0114_
rlabel metal2 69165 22828 69165 22828 0 _0115_
rlabel metal2 57120 16044 57120 16044 0 _0116_
rlabel metal2 68750 22764 68750 22764 0 _0117_
rlabel metal2 68365 22828 68365 22828 0 _0118_
rlabel metal2 67918 22764 67918 22764 0 _0119_
rlabel metal2 67526 22764 67526 22764 0 _0120_
rlabel metal2 67134 22764 67134 22764 0 _0121_
rlabel metal2 66742 22764 66742 22764 0 _0122_
rlabel metal2 66350 22764 66350 22764 0 _0123_
rlabel metal2 65965 22828 65965 22828 0 _0124_
rlabel metal2 65565 22828 65565 22828 0 _0125_
rlabel metal2 65165 22828 65165 22828 0 _0126_
rlabel metal2 57408 16506 57408 16506 0 _0127_
rlabel metal2 22848 19026 22848 19026 0 _0128_
rlabel metal2 26112 18942 26112 18942 0 _0129_
rlabel metal2 29328 18732 29328 18732 0 _0130_
rlabel metal2 32400 19488 32400 19488 0 _0131_
rlabel metal2 35568 20244 35568 20244 0 _0132_
rlabel metal2 38736 20664 38736 20664 0 _0133_
rlabel metal3 41808 20160 41808 20160 0 _0134_
rlabel metal3 40896 17724 40896 17724 0 _0135_
rlabel metal3 40944 13440 40944 13440 0 _0136_
rlabel metal2 39840 14784 39840 14784 0 _0137_
rlabel metal2 37344 15456 37344 15456 0 _0138_
rlabel metal2 31008 15918 31008 15918 0 _0139_
rlabel metal2 33024 13734 33024 13734 0 _0140_
rlabel metal3 34368 11928 34368 11928 0 _0141_
rlabel metal2 36384 10458 36384 10458 0 _0142_
rlabel metal3 39744 9660 39744 9660 0 _0143_
rlabel metal2 41568 8904 41568 8904 0 _0144_
rlabel metal3 44640 8148 44640 8148 0 _0145_
rlabel metal2 45408 7434 45408 7434 0 _0146_
rlabel metal3 46512 5040 46512 5040 0 _0147_
rlabel metal3 49920 3612 49920 3612 0 _0148_
rlabel metal2 52416 5880 52416 5880 0 _0149_
rlabel metal2 52896 7140 52896 7140 0 _0150_
rlabel metal3 51504 9660 51504 9660 0 _0151_
rlabel metal3 49488 11088 49488 11088 0 _0152_
rlabel metal3 46896 11928 46896 11928 0 _0153_
rlabel metal2 46848 11970 46848 11970 0 _0154_
rlabel metal2 45984 15792 45984 15792 0 _0155_
rlabel metal2 46992 18312 46992 18312 0 _0156_
rlabel metal3 49056 16212 49056 16212 0 _0157_
rlabel metal3 51072 14196 51072 14196 0 _0158_
rlabel metal2 54720 13734 54720 13734 0 _0159_
rlabel metal3 55776 13020 55776 13020 0 _0160_
rlabel metal3 57264 10416 57264 10416 0 _0161_
rlabel metal2 55968 8316 55968 8316 0 _0162_
rlabel metal3 57456 6300 57456 6300 0 _0163_
rlabel metal2 58848 5250 58848 5250 0 _0164_
rlabel metal3 56640 3528 56640 3528 0 _0165_
rlabel metal2 53472 1848 53472 1848 0 _0166_
rlabel metal3 59088 1344 59088 1344 0 _0167_
rlabel metal3 62160 1344 62160 1344 0 _0168_
rlabel metal2 62880 3822 62880 3822 0 _0169_
rlabel metal2 62976 5250 62976 5250 0 _0170_
rlabel metal2 62208 7434 62208 7434 0 _0171_
rlabel metal3 63552 9576 63552 9576 0 _0172_
rlabel metal2 63648 11676 63648 11676 0 _0173_
rlabel metal2 61344 12684 61344 12684 0 _0174_
rlabel metal2 64656 13440 64656 13440 0 _0175_
rlabel metal2 68256 14364 68256 14364 0 _0176_
rlabel metal3 68208 11592 68208 11592 0 _0177_
rlabel metal2 66912 9828 66912 9828 0 _0178_
rlabel metal2 68736 8064 68736 8064 0 _0179_
rlabel metal3 69504 5880 69504 5880 0 _0180_
rlabel metal2 66048 1134 66048 1134 0 _0181_
rlabel metal3 69168 3612 69168 3612 0 _0182_
rlabel metal2 71376 2016 71376 2016 0 _0183_
rlabel metal2 75648 1848 75648 1848 0 _0184_
rlabel metal2 74496 4158 74496 4158 0 _0185_
rlabel metal2 76032 5502 76032 5502 0 _0186_
rlabel metal2 75552 7686 75552 7686 0 _0187_
rlabel metal2 75984 9324 75984 9324 0 _0188_
rlabel metal2 72480 11382 72480 11382 0 _0189_
rlabel metal2 74400 13020 74400 13020 0 _0190_
rlabel metal2 72192 14322 72192 14322 0 _0191_
rlabel metal2 73248 25620 73248 25620 0 _0192_
rlabel metal2 74880 27132 74880 27132 0 _0193_
rlabel metal2 75360 28392 75360 28392 0 _0194_
rlabel metal3 74544 30828 74544 30828 0 _0195_
rlabel metal3 75408 33432 75408 33432 0 _0196_
rlabel metal2 76128 34734 76128 34734 0 _0197_
rlabel metal2 76224 36918 76224 36918 0 _0198_
rlabel metal2 73824 37002 73824 37002 0 _0199_
rlabel metal2 71328 34440 71328 34440 0 _0200_
rlabel metal2 65760 36582 65760 36582 0 _0201_
rlabel metal3 65568 35784 65568 35784 0 _0202_
rlabel metal2 66384 33684 66384 33684 0 _0203_
rlabel metal3 69648 32340 69648 32340 0 _0204_
rlabel metal3 69600 29736 69600 29736 0 _0205_
rlabel metal2 67680 29442 67680 29442 0 _0206_
rlabel metal2 69216 27216 69216 27216 0 _0207_
rlabel metal2 67776 26418 67776 26418 0 _0208_
rlabel metal3 63216 26208 63216 26208 0 _0209_
rlabel metal2 61920 28014 61920 28014 0 _0210_
rlabel metal2 63168 30534 63168 30534 0 _0211_
rlabel metal3 61536 31248 61536 31248 0 _0212_
rlabel metal3 60864 34524 60864 34524 0 _0213_
rlabel metal2 62016 37086 62016 37086 0 _0214_
rlabel metal2 55968 37674 55968 37674 0 _0215_
rlabel metal3 55008 36792 55008 36792 0 _0216_
rlabel metal2 57984 34440 57984 34440 0 _0217_
rlabel metal3 58752 30744 58752 30744 0 _0218_
rlabel metal3 58656 27720 58656 27720 0 _0219_
rlabel metal2 57504 25620 57504 25620 0 _0220_
rlabel metal2 56544 26292 56544 26292 0 _0221_
rlabel metal2 54576 27468 54576 27468 0 _0222_
rlabel metal2 52800 30870 52800 30870 0 _0223_
rlabel metal2 54048 33978 54048 33978 0 _0224_
rlabel metal2 50928 34608 50928 34608 0 _0225_
rlabel metal2 46176 34650 46176 34650 0 _0226_
rlabel metal2 48912 33432 48912 33432 0 _0227_
rlabel metal2 48096 30954 48096 30954 0 _0228_
rlabel metal2 48864 27930 48864 27930 0 _0229_
rlabel metal3 50208 26208 50208 26208 0 _0230_
rlabel metal2 48000 23646 48000 23646 0 _0231_
rlabel metal2 47712 21042 47712 21042 0 _0232_
rlabel metal2 45216 21882 45216 21882 0 _0233_
rlabel metal2 44448 24318 44448 24318 0 _0234_
rlabel metal2 44064 25578 44064 25578 0 _0235_
rlabel metal2 45984 27930 45984 27930 0 _0236_
rlabel metal3 44352 28980 44352 28980 0 _0237_
rlabel metal3 41472 30408 41472 30408 0 _0238_
rlabel metal3 39792 28560 39792 28560 0 _0239_
rlabel metal3 39168 27720 39168 27720 0 _0240_
rlabel metal2 37248 25578 37248 25578 0 _0241_
rlabel metal3 38784 22512 38784 22512 0 _0242_
rlabel metal3 35520 24024 35520 24024 0 _0243_
rlabel metal2 34752 25830 34752 25830 0 _0244_
rlabel metal3 31200 24696 31200 24696 0 _0245_
rlabel metal3 29520 23184 29520 23184 0 _0246_
rlabel metal2 28272 20748 28272 20748 0 _0247_
rlabel metal2 8400 18648 8400 18648 0 _0248_
rlabel metal2 2976 3738 2976 3738 0 _0249_
rlabel metal2 2208 5334 2208 5334 0 _0250_
rlabel metal3 1872 6636 1872 6636 0 _0251_
rlabel metal3 1776 8148 1776 8148 0 _0252_
rlabel metal3 1920 10332 1920 10332 0 _0253_
rlabel metal2 2112 13272 2112 13272 0 _0254_
rlabel metal3 1536 14952 1536 14952 0 _0255_
rlabel metal3 22944 17640 22944 17640 0 _0256_
rlabel metal2 27072 17220 27072 17220 0 _0257_
rlabel metal3 30240 17640 30240 17640 0 _0258_
rlabel metal2 32640 18522 32640 18522 0 _0259_
rlabel metal3 36000 18648 36000 18648 0 _0260_
rlabel metal2 38784 18858 38784 18858 0 _0261_
rlabel metal2 44064 18942 44064 18942 0 _0262_
rlabel metal3 43008 17640 43008 17640 0 _0263_
rlabel metal2 43056 13188 43056 13188 0 _0264_
rlabel metal2 40368 15708 40368 15708 0 _0265_
rlabel metal3 37680 16464 37680 16464 0 _0266_
rlabel metal2 33888 17010 33888 17010 0 _0267_
rlabel metal2 31440 13860 31440 13860 0 _0268_
rlabel metal2 36912 11928 36912 11928 0 _0269_
rlabel metal2 39216 11928 39216 11928 0 _0270_
rlabel metal2 42336 11760 42336 11760 0 _0271_
rlabel metal2 44160 10920 44160 10920 0 _0272_
rlabel metal3 46560 10080 46560 10080 0 _0273_
rlabel metal2 48768 7476 48768 7476 0 _0274_
rlabel metal2 48912 5880 48912 5880 0 _0275_
rlabel metal2 52320 4242 52320 4242 0 _0276_
rlabel metal3 54432 6552 54432 6552 0 _0277_
rlabel metal2 54144 7938 54144 7938 0 _0278_
rlabel metal3 53616 10752 53616 10752 0 _0279_
rlabel metal2 51840 11844 51840 11844 0 _0280_
rlabel metal3 49296 13104 49296 13104 0 _0281_
rlabel metal2 47712 13986 47712 13986 0 _0282_
rlabel metal2 45984 16506 45984 16506 0 _0283_
rlabel metal3 49392 19152 49392 19152 0 _0284_
rlabel metal2 50304 17808 50304 17808 0 _0285_
rlabel metal2 53184 15666 53184 15666 0 _0286_
rlabel metal2 56928 15246 56928 15246 0 _0287_
rlabel metal2 58752 13482 58752 13482 0 _0288_
rlabel metal3 59136 11592 59136 11592 0 _0289_
rlabel metal2 59232 8694 59232 8694 0 _0290_
rlabel metal2 60768 7518 60768 7518 0 _0291_
rlabel metal2 61248 5922 61248 5922 0 _0292_
rlabel metal2 55920 5124 55920 5124 0 _0293_
rlabel metal2 56640 2226 56640 2226 0 _0294_
rlabel metal3 59280 3444 59280 3444 0 _0295_
rlabel metal2 64512 2058 64512 2058 0 _0296_
rlabel metal2 66240 3822 66240 3822 0 _0297_
rlabel metal2 66480 5880 66480 5880 0 _0298_
rlabel metal2 65808 8148 65808 8148 0 _0299_
rlabel metal2 65280 10458 65280 10458 0 _0300_
rlabel metal2 64704 11928 64704 11928 0 _0301_
rlabel metal2 60864 14952 60864 14952 0 _0302_
rlabel metal2 65424 14952 65424 14952 0 _0303_
rlabel metal2 70368 14994 70368 14994 0 _0304_
rlabel metal2 70464 12432 70464 12432 0 _0305_
rlabel metal3 70176 9324 70176 9324 0 _0306_
rlabel metal2 71520 8358 71520 8358 0 _0307_
rlabel metal2 72000 6678 72000 6678 0 _0308_
rlabel metal2 68880 1344 68880 1344 0 _0309_
rlabel metal2 71904 4410 71904 4410 0 _0310_
rlabel metal2 74016 1386 74016 1386 0 _0311_
rlabel metal2 79488 1176 79488 1176 0 _0312_
rlabel metal2 77088 4410 77088 4410 0 _0313_
rlabel metal2 77136 5880 77136 5880 0 _0314_
rlabel metal2 77088 8358 77088 8358 0 _0315_
rlabel metal2 77136 9660 77136 9660 0 _0316_
rlabel metal2 76416 12222 76416 12222 0 _0317_
rlabel metal2 76512 13734 76512 13734 0 _0318_
rlabel metal2 76224 14784 76224 14784 0 _0319_
rlabel metal3 76512 25200 76512 25200 0 _0320_
rlabel metal3 76992 26292 76992 26292 0 _0321_
rlabel metal2 76800 28602 76800 28602 0 _0322_
rlabel metal2 77088 30366 77088 30366 0 _0323_
rlabel metal2 77184 32256 77184 32256 0 _0324_
rlabel metal2 77424 34524 77424 34524 0 _0325_
rlabel metal3 76848 36540 76848 36540 0 _0326_
rlabel metal2 73344 37086 73344 37086 0 _0327_
rlabel metal2 72192 34440 72192 34440 0 _0328_
rlabel metal2 69024 37704 69024 37704 0 _0329_
rlabel metal2 67008 34650 67008 34650 0 _0330_
rlabel metal2 66480 31584 66480 31584 0 _0331_
rlabel metal2 72096 32844 72096 32844 0 _0332_
rlabel metal2 71664 30072 71664 30072 0 _0333_
rlabel metal2 71280 27804 71280 27804 0 _0334_
rlabel metal2 70752 24780 70752 24780 0 _0335_
rlabel metal2 67776 24990 67776 24990 0 _0336_
rlabel metal2 64032 24990 64032 24990 0 _0337_
rlabel metal2 65136 27468 65136 27468 0 _0338_
rlabel metal2 65760 29106 65760 29106 0 _0339_
rlabel metal2 63024 31584 63024 31584 0 _0340_
rlabel metal3 62880 34272 62880 34272 0 _0341_
rlabel metal3 63936 37968 63936 37968 0 _0342_
rlabel metal2 59184 36876 59184 36876 0 _0343_
rlabel metal3 55392 35364 55392 35364 0 _0344_
rlabel metal3 58560 32760 58560 32760 0 _0345_
rlabel metal2 60576 29316 60576 29316 0 _0346_
rlabel metal2 60432 27720 60432 27720 0 _0347_
rlabel metal2 60144 25284 60144 25284 0 _0348_
rlabel metal2 55392 24318 55392 24318 0 _0349_
rlabel metal2 56208 28560 56208 28560 0 _0350_
rlabel metal2 56112 30828 56112 30828 0 _0351_
rlabel metal2 55680 32928 55680 32928 0 _0352_
rlabel metal2 52272 34944 52272 34944 0 _0353_
rlabel metal2 45840 32256 45840 32256 0 _0354_
rlabel metal2 51072 31584 51072 31584 0 _0355_
rlabel metal2 51168 29316 51168 29316 0 _0356_
rlabel metal3 51840 27720 51840 27720 0 _0357_
rlabel metal2 52080 24444 52080 24444 0 _0358_
rlabel metal2 51744 23856 51744 23856 0 _0359_
rlabel metal2 50352 20748 50352 20748 0 _0360_
rlabel metal2 45744 20580 45744 20580 0 _0361_
rlabel metal2 46320 22848 46320 22848 0 _0362_
rlabel metal2 47184 24444 47184 24444 0 _0363_
rlabel metal2 47136 27090 47136 27090 0 _0364_
rlabel metal2 46560 30114 46560 30114 0 _0365_
rlabel metal2 43968 31626 43968 31626 0 _0366_
rlabel metal2 41952 28392 41952 28392 0 _0367_
rlabel metal2 41664 26292 41664 26292 0 _0368_
rlabel metal3 40656 23688 40656 23688 0 _0369_
rlabel metal2 41088 22134 41088 22134 0 _0370_
rlabel metal3 36048 21756 36048 21756 0 _0371_
rlabel metal2 35712 26502 35712 26502 0 _0372_
rlabel metal2 32976 23268 32976 23268 0 _0373_
rlabel metal2 32544 22092 32544 22092 0 _0374_
rlabel metal3 29040 20664 29040 20664 0 _0375_
rlabel metal2 9312 19320 9312 19320 0 _0376_
rlabel metal2 5280 4200 5280 4200 0 _0377_
rlabel metal3 5712 5880 5712 5880 0 _0378_
rlabel metal2 4896 8148 4896 8148 0 _0379_
rlabel metal3 4656 9576 4656 9576 0 _0380_
rlabel metal2 4992 11760 4992 11760 0 _0381_
rlabel metal3 4848 12684 4848 12684 0 _0382_
rlabel metal2 4608 15708 4608 15708 0 _0383_
rlabel metal2 64416 8694 64416 8694 0 _0384_
rlabel metal2 64128 8820 64128 8820 0 _0385_
rlabel metal2 64128 11424 64128 11424 0 _0386_
rlabel metal2 63264 12432 63264 12432 0 _0387_
rlabel metal3 63504 10416 63504 10416 0 _0388_
rlabel metal2 63072 11802 63072 11802 0 _0389_
rlabel metal2 61056 13734 61056 13734 0 _0390_
rlabel metal2 61152 14448 61152 14448 0 _0391_
rlabel metal2 61632 12432 61632 12432 0 _0392_
rlabel metal3 61584 13020 61584 13020 0 _0393_
rlabel metal2 63936 14784 63936 14784 0 _0394_
rlabel metal3 64512 14700 64512 14700 0 _0395_
rlabel metal2 64320 13482 64320 13482 0 _0396_
rlabel metal3 64224 13020 64224 13020 0 _0397_
rlabel metal2 70320 13188 70320 13188 0 _0398_
rlabel metal2 70176 13482 70176 13482 0 _0399_
rlabel metal2 68064 13944 68064 13944 0 _0400_
rlabel metal2 68352 14217 68352 14217 0 _0401_
rlabel metal3 69696 11928 69696 11928 0 _0402_
rlabel metal3 69600 12516 69600 12516 0 _0403_
rlabel metal2 69216 12348 69216 12348 0 _0404_
rlabel metal4 68928 12348 68928 12348 0 _0405_
rlabel metal2 69936 8652 69936 8652 0 _0406_
rlabel metal2 70080 9912 70080 9912 0 _0407_
rlabel metal2 69024 10458 69024 10458 0 _0408_
rlabel metal2 68256 10206 68256 10206 0 _0409_
rlabel metal2 71520 9198 71520 9198 0 _0410_
rlabel metal3 70176 9240 70176 9240 0 _0411_
rlabel metal2 69024 8736 69024 8736 0 _0412_
rlabel metal2 69600 7896 69600 7896 0 _0413_
rlabel metal2 72192 5670 72192 5670 0 _0414_
rlabel metal3 71136 5544 71136 5544 0 _0415_
rlabel metal2 70080 6300 70080 6300 0 _0416_
rlabel metal2 69696 5628 69696 5628 0 _0417_
rlabel metal2 68640 2184 68640 2184 0 _0418_
rlabel metal2 68736 1008 68736 1008 0 _0419_
rlabel metal2 67680 2406 67680 2406 0 _0420_
rlabel metal2 67392 2184 67392 2184 0 _0421_
rlabel metal2 71184 4956 71184 4956 0 _0422_
rlabel metal3 70272 4704 70272 4704 0 _0423_
rlabel metal2 69120 3360 69120 3360 0 _0424_
rlabel metal2 69552 3444 69552 3444 0 _0425_
rlabel via1 73344 2868 73344 2868 0 _0426_
rlabel metal2 74208 2310 74208 2310 0 _0427_
rlabel metal2 71136 2742 71136 2742 0 _0428_
rlabel metal2 71520 2604 71520 2604 0 _0429_
rlabel metal2 77664 2688 77664 2688 0 _0430_
rlabel metal2 77760 2226 77760 2226 0 _0431_
rlabel metal2 75168 1848 75168 1848 0 _0432_
rlabel metal2 75888 924 75888 924 0 _0433_
rlabel metal2 77280 3360 77280 3360 0 _0434_
rlabel metal2 77376 4242 77376 4242 0 _0435_
rlabel metal2 76368 4032 76368 4032 0 _0436_
rlabel metal2 76128 3654 76128 3654 0 _0437_
rlabel metal2 76992 6720 76992 6720 0 _0438_
rlabel metal2 77328 5628 77328 5628 0 _0439_
rlabel metal2 76128 5208 76128 5208 0 _0440_
rlabel metal2 76176 5628 76176 5628 0 _0441_
rlabel metal2 76848 7980 76848 7980 0 _0442_
rlabel metal2 76704 7434 76704 7434 0 _0443_
rlabel metal2 75840 7098 75840 7098 0 _0444_
rlabel metal2 75600 7140 75600 7140 0 _0445_
rlabel via1 77079 11010 77079 11010 0 _0446_
rlabel metal2 77232 10752 77232 10752 0 _0447_
rlabel metal3 76032 8568 76032 8568 0 _0448_
rlabel metal2 76032 9660 76032 9660 0 _0449_
rlabel metal2 76128 11424 76128 11424 0 _0450_
rlabel metal2 76224 11382 76224 11382 0 _0451_
rlabel metal2 75456 10920 75456 10920 0 _0452_
rlabel metal3 74928 11004 74928 11004 0 _0453_
rlabel metal2 76128 13158 76128 13158 0 _0454_
rlabel metal2 76704 13074 76704 13074 0 _0455_
rlabel metal2 74592 12432 74592 12432 0 _0456_
rlabel metal3 74544 13188 74544 13188 0 _0457_
rlabel metal2 75456 15540 75456 15540 0 _0458_
rlabel metal3 74544 15288 74544 15288 0 _0459_
rlabel metal2 74784 13734 74784 13734 0 _0460_
rlabel metal2 74112 14784 74112 14784 0 _0461_
rlabel via1 76032 25284 76032 25284 0 _0462_
rlabel metal2 76416 25704 76416 25704 0 _0463_
rlabel metal2 74304 24780 74304 24780 0 _0464_
rlabel metal2 74496 26208 74496 26208 0 _0465_
rlabel metal2 76896 27342 76896 27342 0 _0466_
rlabel metal3 75936 27636 75936 27636 0 _0467_
rlabel metal2 75264 26082 75264 26082 0 _0468_
rlabel metal3 75216 26796 75216 26796 0 _0469_
rlabel metal2 76752 29820 76752 29820 0 _0470_
rlabel metal2 76944 28308 76944 28308 0 _0471_
rlabel metal2 75408 27384 75408 27384 0 _0472_
rlabel metal2 75264 28434 75264 28434 0 _0473_
rlabel metal2 76992 30912 76992 30912 0 _0474_
rlabel metal2 77280 30030 77280 30030 0 _0475_
rlabel metal2 75696 30072 75696 30072 0 _0476_
rlabel metal2 75360 30702 75360 30702 0 _0477_
rlabel metal3 78336 32844 78336 32844 0 _0478_
rlabel metal3 77952 33684 77952 33684 0 _0479_
rlabel metal2 75840 32340 75840 32340 0 _0480_
rlabel metal2 76128 33684 76128 33684 0 _0481_
rlabel metal2 77280 35238 77280 35238 0 _0482_
rlabel metal2 77664 34860 77664 34860 0 _0483_
rlabel metal2 76800 34020 76800 34020 0 _0484_
rlabel metal2 76032 35028 76032 35028 0 _0485_
rlabel metal2 77664 36918 77664 36918 0 _0486_
rlabel metal2 76800 36414 76800 36414 0 _0487_
rlabel metal2 76464 36120 76464 36120 0 _0488_
rlabel metal2 75792 36708 75792 36708 0 _0489_
rlabel metal3 73728 35868 73728 35868 0 _0490_
rlabel metal2 73920 37338 73920 37338 0 _0491_
rlabel metal3 74160 37380 74160 37380 0 _0492_
rlabel metal2 73056 37380 73056 37380 0 _0493_
rlabel metal2 72384 35112 72384 35112 0 _0494_
rlabel metal2 72096 34986 72096 34986 0 _0495_
rlabel metal2 72192 35448 72192 35448 0 _0496_
rlabel metal3 71328 35196 71328 35196 0 _0497_
rlabel metal2 68736 37065 68736 37065 0 _0498_
rlabel metal2 68832 37830 68832 37830 0 _0499_
rlabel metal2 69792 36246 69792 36246 0 _0500_
rlabel metal2 68448 38220 68448 38220 0 _0501_
rlabel metal2 67488 35658 67488 35658 0 _0502_
rlabel metal2 67008 35364 67008 35364 0 _0503_
rlabel metal2 67152 35868 67152 35868 0 _0504_
rlabel metal3 66336 35364 66336 35364 0 _0505_
rlabel metal2 65664 32172 65664 32172 0 _0506_
rlabel metal2 66624 31668 66624 31668 0 _0507_
rlabel metal3 66528 34188 66528 34188 0 _0508_
rlabel metal2 66432 32844 66432 32844 0 _0509_
rlabel metal2 72384 32172 72384 32172 0 _0510_
rlabel metal2 72144 33684 72144 33684 0 _0511_
rlabel metal2 69792 32424 69792 32424 0 _0512_
rlabel metal2 70176 32172 70176 32172 0 _0513_
rlabel metal2 71616 30912 71616 30912 0 _0514_
rlabel metal2 71712 29736 71712 29736 0 _0515_
rlabel metal2 71136 30324 71136 30324 0 _0516_
rlabel metal2 70848 30492 70848 30492 0 _0517_
rlabel metal2 70896 27636 70896 27636 0 _0518_
rlabel metal2 70752 28140 70752 28140 0 _0519_
rlabel metal2 70176 29904 70176 29904 0 _0520_
rlabel metal2 70080 29316 70080 29316 0 _0521_
rlabel metal2 71808 25998 71808 25998 0 _0522_
rlabel metal2 71904 26628 71904 26628 0 _0523_
rlabel metal2 69888 27552 69888 27552 0 _0524_
rlabel metal2 69648 26292 69648 26292 0 _0525_
rlabel metal2 68352 25830 68352 25830 0 _0526_
rlabel metal2 67872 25914 67872 25914 0 _0527_
rlabel metal2 67968 26250 67968 26250 0 _0528_
rlabel metal2 67584 26124 67584 26124 0 _0529_
rlabel metal2 63792 24612 63792 24612 0 _0530_
rlabel metal2 64128 24864 64128 24864 0 _0531_
rlabel metal2 64992 26040 64992 26040 0 _0532_
rlabel metal2 64608 26124 64608 26124 0 _0533_
rlabel metal2 64800 27846 64800 27846 0 _0534_
rlabel metal3 64368 27636 64368 27636 0 _0535_
rlabel metal2 63792 27048 63792 27048 0 _0536_
rlabel metal2 64080 27636 64080 27636 0 _0537_
rlabel metal2 64992 29820 64992 29820 0 _0538_
rlabel metal2 64800 29442 64800 29442 0 _0539_
rlabel metal3 63744 29316 63744 29316 0 _0540_
rlabel metal2 63648 29820 63648 29820 0 _0541_
rlabel metal2 63936 32088 63936 32088 0 _0542_
rlabel metal2 63264 31458 63264 31458 0 _0543_
rlabel metal2 62832 30828 62832 30828 0 _0544_
rlabel metal2 62592 32004 62592 32004 0 _0545_
rlabel metal2 62688 33768 62688 33768 0 _0546_
rlabel metal2 62784 34062 62784 34062 0 _0547_
rlabel metal2 62304 34062 62304 34062 0 _0548_
rlabel metal2 61872 34356 61872 34356 0 _0549_
rlabel metal3 63936 36708 63936 36708 0 _0550_
rlabel metal2 63744 37380 63744 37380 0 _0551_
rlabel metal2 61440 35910 61440 35910 0 _0552_
rlabel metal2 61824 36708 61824 36708 0 _0553_
rlabel metal2 58848 36162 58848 36162 0 _0554_
rlabel metal2 59328 36792 59328 36792 0 _0555_
rlabel metal2 60288 37170 60288 37170 0 _0556_
rlabel metal3 58512 37212 58512 37212 0 _0557_
rlabel metal2 54912 35028 54912 35028 0 _0558_
rlabel metal2 55296 35238 55296 35238 0 _0559_
rlabel metal3 56448 36876 56448 36876 0 _0560_
rlabel metal2 55776 35952 55776 35952 0 _0561_
rlabel metal2 59232 32088 59232 32088 0 _0562_
rlabel metal3 57696 33768 57696 33768 0 _0563_
rlabel metal2 57504 34650 57504 34650 0 _0564_
rlabel metal2 58368 33894 58368 33894 0 _0565_
rlabel metal2 60864 29316 60864 29316 0 _0566_
rlabel metal2 60960 29736 60960 29736 0 _0567_
rlabel metal2 59904 31626 59904 31626 0 _0568_
rlabel metal2 59232 30576 59232 30576 0 _0569_
rlabel metal2 60672 27888 60672 27888 0 _0570_
rlabel metal3 60576 28308 60576 28308 0 _0571_
rlabel metal2 60192 27888 60192 27888 0 _0572_
rlabel metal2 59664 27636 59664 27636 0 _0573_
rlabel metal2 59520 25998 59520 25998 0 _0574_
rlabel metal2 59808 26040 59808 26040 0 _0575_
rlabel metal3 58800 26124 58800 26124 0 _0576_
rlabel metal2 58320 24780 58320 24780 0 _0577_
rlabel metal2 55200 26040 55200 26040 0 _0578_
rlabel metal3 55824 25956 55824 25956 0 _0579_
rlabel metal2 56640 26040 56640 26040 0 _0580_
rlabel metal2 56352 26460 56352 26460 0 _0581_
rlabel metal2 55872 29190 55872 29190 0 _0582_
rlabel metal2 56448 27972 56448 27972 0 _0583_
rlabel metal2 54912 27468 54912 27468 0 _0584_
rlabel metal2 54672 27636 54672 27636 0 _0585_
rlabel metal2 55776 30912 55776 30912 0 _0586_
rlabel metal3 55440 30660 55440 30660 0 _0587_
rlabel metal2 54816 30366 54816 30366 0 _0588_
rlabel metal2 54576 30660 54576 30660 0 _0589_
rlabel metal2 55296 34356 55296 34356 0 _0590_
rlabel metal2 55104 34062 55104 34062 0 _0591_
rlabel metal2 54240 33348 54240 33348 0 _0592_
rlabel metal2 53952 33600 53952 33600 0 _0593_
rlabel metal2 51264 35448 51264 35448 0 _0594_
rlabel metal2 52128 35147 52128 35147 0 _0595_
rlabel metal2 51264 34440 51264 34440 0 _0596_
rlabel metal2 50880 34356 50880 34356 0 _0597_
rlabel metal3 47328 32844 47328 32844 0 _0598_
rlabel metal2 46800 34188 46800 34188 0 _0599_
rlabel metal3 48048 34524 48048 34524 0 _0600_
rlabel metal2 46560 33852 46560 33852 0 _0601_
rlabel metal2 51072 32550 51072 32550 0 _0602_
rlabel metal3 50064 33684 50064 33684 0 _0603_
rlabel metal2 48864 31668 48864 31668 0 _0604_
rlabel metal2 48864 33684 48864 33684 0 _0605_
rlabel metal2 50976 30366 50976 30366 0 _0606_
rlabel metal2 50880 30786 50880 30786 0 _0607_
rlabel metal2 49536 31416 49536 31416 0 _0608_
rlabel metal3 49488 29820 49488 29820 0 _0609_
rlabel metal2 51888 28308 51888 28308 0 _0610_
rlabel metal3 50976 28476 50976 28476 0 _0611_
rlabel metal2 50304 28602 50304 28602 0 _0612_
rlabel metal3 50256 28308 50256 28308 0 _0613_
rlabel metal2 51360 25284 51360 25284 0 _0614_
rlabel metal2 51168 24906 51168 24906 0 _0615_
rlabel metal3 51216 26124 51216 26124 0 _0616_
rlabel metal2 50880 25704 50880 25704 0 _0617_
rlabel metal2 50976 22986 50976 22986 0 _0618_
rlabel metal2 51264 23478 51264 23478 0 _0619_
rlabel metal2 50880 24066 50880 24066 0 _0620_
rlabel metal2 50016 23520 50016 23520 0 _0621_
rlabel metal2 49728 21504 49728 21504 0 _0622_
rlabel metal3 50304 21588 50304 21588 0 _0623_
rlabel metal2 49248 21588 49248 21588 0 _0624_
rlabel metal2 48864 21840 48864 21840 0 _0625_
rlabel metal2 45984 21042 45984 21042 0 _0626_
rlabel metal2 46080 21504 46080 21504 0 _0627_
rlabel metal2 46320 21000 46320 21000 0 _0628_
rlabel metal2 45120 21504 45120 21504 0 _0629_
rlabel metal2 45888 23772 45888 23772 0 _0630_
rlabel metal3 45360 23772 45360 23772 0 _0631_
rlabel metal2 44736 23520 44736 23520 0 _0632_
rlabel metal3 44208 23772 44208 23772 0 _0633_
rlabel via1 46271 25284 46271 25284 0 _0634_
rlabel metal3 45312 25452 45312 25452 0 _0635_
rlabel metal2 45024 25032 45024 25032 0 _0636_
rlabel metal2 44352 25116 44352 25116 0 _0637_
rlabel metal2 46848 27888 46848 27888 0 _0638_
rlabel metal3 47040 28224 47040 28224 0 _0639_
rlabel metal2 46512 26292 46512 26292 0 _0640_
rlabel metal2 45504 28308 45504 28308 0 _0641_
rlabel metal2 45888 29820 45888 29820 0 _0642_
rlabel metal3 45648 30408 45648 30408 0 _0643_
rlabel metal3 45024 28560 45024 28560 0 _0644_
rlabel metal2 45168 29148 45168 29148 0 _0645_
rlabel metal2 42912 31920 42912 31920 0 _0646_
rlabel metal2 42960 30660 42960 30660 0 _0647_
rlabel metal2 43104 30576 43104 30576 0 _0648_
rlabel metal2 42816 30612 42816 30612 0 _0649_
rlabel metal2 41232 29820 41232 29820 0 _0650_
rlabel metal2 42144 29442 42144 29442 0 _0651_
rlabel metal2 41376 28602 41376 28602 0 _0652_
rlabel metal2 41040 28308 41040 28308 0 _0653_
rlabel metal2 41280 27342 41280 27342 0 _0654_
rlabel metal2 41136 27384 41136 27384 0 _0655_
rlabel metal2 40752 27636 40752 27636 0 _0656_
rlabel metal2 40272 26796 40272 26796 0 _0657_
rlabel metal2 40272 25284 40272 25284 0 _0658_
rlabel metal2 40368 25536 40368 25536 0 _0659_
rlabel metal2 39552 26040 39552 26040 0 _0660_
rlabel metal2 40128 25452 40128 25452 0 _0661_
rlabel metal2 41088 23583 41088 23583 0 _0662_
rlabel metal3 40032 22260 40032 22260 0 _0663_
rlabel metal2 39456 22260 39456 22260 0 _0664_
rlabel metal2 39024 22260 39024 22260 0 _0665_
rlabel metal3 37056 23268 37056 23268 0 _0666_
rlabel metal2 36336 23352 36336 23352 0 _0667_
rlabel metal2 37920 23310 37920 23310 0 _0668_
rlabel metal2 35712 23520 35712 23520 0 _0669_
rlabel metal2 35232 26376 35232 26376 0 _0670_
rlabel metal2 35616 26544 35616 26544 0 _0671_
rlabel metal2 35040 25410 35040 25410 0 _0672_
rlabel metal2 34656 25284 34656 25284 0 _0673_
rlabel metal2 32544 23520 32544 23520 0 _0674_
rlabel metal2 32448 23352 32448 23352 0 _0675_
rlabel metal2 33312 24864 33312 24864 0 _0676_
rlabel metal2 32352 24612 32352 24612 0 _0677_
rlabel metal2 31680 22008 31680 22008 0 _0678_
rlabel metal3 32064 22344 32064 22344 0 _0679_
rlabel metal3 31152 23268 31152 23268 0 _0680_
rlabel metal2 30672 22260 30672 22260 0 _0681_
rlabel metal2 28704 20076 28704 20076 0 _0682_
rlabel metal3 28704 20748 28704 20748 0 _0683_
rlabel metal2 28704 21588 28704 21588 0 _0684_
rlabel metal2 28224 21588 28224 21588 0 _0685_
rlabel metal2 8544 17808 8544 17808 0 _0686_
rlabel metal2 8544 19026 8544 19026 0 _0687_
rlabel metal2 26688 19488 26688 19488 0 _0688_
rlabel metal2 8832 18774 8832 18774 0 _0689_
rlabel metal2 4272 3444 4272 3444 0 _0690_
rlabel metal3 3984 4116 3984 4116 0 _0691_
rlabel metal2 3024 2856 3024 2856 0 _0692_
rlabel metal2 2832 2604 2832 2604 0 _0693_
rlabel metal2 3696 4956 3696 4956 0 _0694_
rlabel metal2 2304 5040 2304 5040 0 _0695_
rlabel metal2 2400 4662 2400 4662 0 _0696_
rlabel metal2 2016 4956 2016 4956 0 _0697_
rlabel metal2 4176 7140 4176 7140 0 _0698_
rlabel metal2 2304 6762 2304 6762 0 _0699_
rlabel metal2 2400 6384 2400 6384 0 _0700_
rlabel metal2 2112 7224 2112 7224 0 _0701_
rlabel metal2 3744 9450 3744 9450 0 _0702_
rlabel metal2 2496 8232 2496 8232 0 _0703_
rlabel metal2 2592 7896 2592 7896 0 _0704_
rlabel metal2 2304 8736 2304 8736 0 _0705_
rlabel metal2 4128 11424 4128 11424 0 _0706_
rlabel metal2 4224 10458 4224 10458 0 _0707_
rlabel metal2 2496 10248 2496 10248 0 _0708_
rlabel metal2 2256 10164 2256 10164 0 _0709_
rlabel metal2 6624 13482 6624 13482 0 _0710_
rlabel metal3 2304 13188 2304 13188 0 _0711_
rlabel metal2 2352 12348 2352 12348 0 _0712_
rlabel metal2 1920 12936 1920 12936 0 _0713_
rlabel metal2 3360 15876 3360 15876 0 _0714_
rlabel metal2 2208 15204 2208 15204 0 _0715_
rlabel metal2 2304 14448 2304 14448 0 _0716_
rlabel metal2 1920 14700 1920 14700 0 _0717_
rlabel metal2 22944 17502 22944 17502 0 _0718_
rlabel metal3 27648 16128 27648 16128 0 _0719_
rlabel metal2 30240 17502 30240 17502 0 _0720_
rlabel metal2 33360 17976 33360 17976 0 _0721_
rlabel metal2 36480 18018 36480 18018 0 _0722_
rlabel metal2 38592 19320 38592 19320 0 _0723_
rlabel metal3 44400 18564 44400 18564 0 _0724_
rlabel metal2 43008 17094 43008 17094 0 _0725_
rlabel metal3 43248 14700 43248 14700 0 _0726_
rlabel metal2 40752 15540 40752 15540 0 _0727_
rlabel metal2 37728 16506 37728 16506 0 _0728_
rlabel metal2 34080 17178 34080 17178 0 _0729_
rlabel metal2 31776 14658 31776 14658 0 _0730_
rlabel metal2 36672 13032 36672 13032 0 _0731_
rlabel metal2 39072 10248 39072 10248 0 _0732_
rlabel metal2 41856 11970 41856 11970 0 _0733_
rlabel metal2 43680 10920 43680 10920 0 _0734_
rlabel metal2 46560 10290 46560 10290 0 _0735_
rlabel metal3 49488 8652 49488 8652 0 _0736_
rlabel metal3 48912 5040 48912 5040 0 _0737_
rlabel metal2 51840 4998 51840 4998 0 _0738_
rlabel metal2 54816 6090 54816 6090 0 _0739_
rlabel metal2 54336 8610 54336 8610 0 _0740_
rlabel metal2 53664 11130 53664 11130 0 _0741_
rlabel metal2 51648 11970 51648 11970 0 _0742_
rlabel metal3 49488 12516 49488 12516 0 _0743_
rlabel metal2 47904 14658 47904 14658 0 _0744_
rlabel metal4 46272 17304 46272 17304 0 _0745_
rlabel metal2 49440 18690 49440 18690 0 _0746_
rlabel metal3 50640 17136 50640 17136 0 _0747_
rlabel metal2 52896 16296 52896 16296 0 _0748_
rlabel metal2 57216 14784 57216 14784 0 _0749_
rlabel metal2 59040 13482 59040 13482 0 _0750_
rlabel metal2 59136 11970 59136 11970 0 _0751_
rlabel metal3 59760 8652 59760 8652 0 _0752_
rlabel metal2 60576 7434 60576 7434 0 _0753_
rlabel metal2 61920 5754 61920 5754 0 _0754_
rlabel metal3 56160 4956 56160 4956 0 _0755_
rlabel metal2 57024 1260 57024 1260 0 _0756_
rlabel metal2 59280 3192 59280 3192 0 _0757_
rlabel metal2 64512 2646 64512 2646 0 _0758_
rlabel metal2 66480 3444 66480 3444 0 _0759_
rlabel metal2 66672 5628 66672 5628 0 _0760_
rlabel metal2 65904 7392 65904 7392 0 _0761_
rlabel metal2 65376 10290 65376 10290 0 _0762_
rlabel metal2 64320 11970 64320 11970 0 _0763_
rlabel metal3 61776 14700 61776 14700 0 _0764_
rlabel metal2 65088 14994 65088 14994 0 _0765_
rlabel metal2 71040 14280 71040 14280 0 _0766_
rlabel metal2 70560 11970 70560 11970 0 _0767_
rlabel metal3 70512 9492 70512 9492 0 _0768_
rlabel metal2 71760 7980 71760 7980 0 _0769_
rlabel metal2 72672 6510 72672 6510 0 _0770_
rlabel metal2 68640 1344 68640 1344 0 _0771_
rlabel metal2 72192 4242 72192 4242 0 _0772_
rlabel metal2 74352 1932 74352 1932 0 _0773_
rlabel metal2 78528 1848 78528 1848 0 _0774_
rlabel metal2 77760 4242 77760 4242 0 _0775_
rlabel metal2 77520 5628 77520 5628 0 _0776_
rlabel metal3 77664 7980 77664 7980 0 _0777_
rlabel metal2 77376 9408 77376 9408 0 _0778_
rlabel metal2 76752 11676 76752 11676 0 _0779_
rlabel metal2 76800 13272 76800 13272 0 _0780_
rlabel metal2 75936 14406 75936 14406 0 _0781_
rlabel metal2 76608 24738 76608 24738 0 _0782_
rlabel metal2 77184 26124 77184 26124 0 _0783_
rlabel metal2 77088 28224 77088 28224 0 _0784_
rlabel metal2 77376 30156 77376 30156 0 _0785_
rlabel metal3 77184 33432 77184 33432 0 _0786_
rlabel metal2 77760 34440 77760 34440 0 _0787_
rlabel metal3 77568 36708 77568 36708 0 _0788_
rlabel metal2 73728 36582 73728 36582 0 _0789_
rlabel metal2 71712 34062 71712 34062 0 _0790_
rlabel metal3 69072 37800 69072 37800 0 _0791_
rlabel metal3 67440 34356 67440 34356 0 _0792_
rlabel metal2 66720 31290 66720 31290 0 _0793_
rlabel metal2 72288 33642 72288 33642 0 _0794_
rlabel metal3 71952 29820 71952 29820 0 _0795_
rlabel metal2 71328 27510 71328 27510 0 _0796_
rlabel metal3 71376 24612 71376 24612 0 _0797_
rlabel metal2 67968 24696 67968 24696 0 _0798_
rlabel metal2 64224 24696 64224 24696 0 _0799_
rlabel metal2 65472 27594 65472 27594 0 _0800_
rlabel metal2 65952 29778 65952 29778 0 _0801_
rlabel metal2 63378 31379 63378 31379 0 _0802_
rlabel metal2 63168 33894 63168 33894 0 _0803_
rlabel metal2 63840 38304 63840 38304 0 _0804_
rlabel metal2 59424 36792 59424 36792 0 _0805_
rlabel via1 55410 35190 55410 35190 0 _0806_
rlabel metal3 58752 33432 58752 33432 0 _0807_
rlabel metal3 60960 29148 60960 29148 0 _0808_
rlabel metal2 60864 27552 60864 27552 0 _0809_
rlabel metal2 60192 24780 60192 24780 0 _0810_
rlabel metal2 55680 24108 55680 24108 0 _0811_
rlabel metal2 56544 28224 56544 28224 0 _0812_
rlabel metal2 56256 30618 56256 30618 0 _0813_
rlabel metal3 55056 32844 55056 32844 0 _0814_
rlabel metal2 51840 34524 51840 34524 0 _0815_
rlabel metal2 45984 32802 45984 32802 0 _0816_
rlabel metal2 51504 31332 51504 31332 0 _0817_
rlabel metal2 50832 29148 50832 29148 0 _0818_
rlabel metal2 52128 27132 52128 27132 0 _0819_
rlabel metal2 52416 24696 52416 24696 0 _0820_
rlabel metal2 51648 23520 51648 23520 0 _0821_
rlabel metal2 50880 21882 50880 21882 0 _0822_
rlabel metal2 45792 21126 45792 21126 0 _0823_
rlabel metal3 45744 23100 45744 23100 0 _0824_
rlabel metal2 47472 24612 47472 24612 0 _0825_
rlabel metal2 47424 27678 47424 27678 0 _0826_
rlabel metal2 46272 30366 46272 30366 0 _0827_
rlabel metal2 43392 30786 43392 30786 0 _0828_
rlabel metal2 41664 28854 41664 28854 0 _0829_
rlabel metal2 41376 26250 41376 26250 0 _0830_
rlabel metal3 40848 24612 40848 24612 0 _0831_
rlabel metal2 41184 22008 41184 22008 0 _0832_
rlabel metal2 36480 21504 36480 21504 0 _0833_
rlabel metal2 35472 25536 35472 25536 0 _0834_
rlabel metal3 33168 23100 33168 23100 0 _0835_
rlabel metal2 32160 21966 32160 21966 0 _0836_
rlabel metal2 28992 21042 28992 21042 0 _0837_
rlabel metal2 9504 18942 9504 18942 0 _0838_
rlabel metal2 4800 4158 4800 4158 0 _0839_
rlabel metal2 3936 5082 3936 5082 0 _0840_
rlabel metal2 4992 7392 4992 7392 0 _0841_
rlabel metal2 4896 9030 4896 9030 0 _0842_
rlabel metal2 4992 11214 4992 11214 0 _0843_
rlabel metal3 4992 14616 4992 14616 0 _0844_
rlabel metal3 4512 15540 4512 15540 0 _0845_
rlabel metal2 3840 29190 3840 29190 0 _0846_
rlabel metal3 7296 19992 7296 19992 0 _0847_
rlabel metal2 23424 17796 23424 17796 0 _0848_
rlabel metal2 22848 18102 22848 18102 0 _0849_
rlabel metal2 1920 22596 1920 22596 0 _0850_
rlabel metal2 1920 20076 1920 20076 0 _0851_
rlabel metal2 22272 20454 22272 20454 0 _0852_
rlabel via1 22656 19229 22656 19229 0 _0853_
rlabel metal2 26592 17808 26592 17808 0 _0854_
rlabel metal2 26304 17976 26304 17976 0 _0855_
rlabel metal2 25920 18480 25920 18480 0 _0856_
rlabel metal2 26304 18564 26304 18564 0 _0857_
rlabel metal2 31104 18480 31104 18480 0 _0858_
rlabel metal2 30144 18018 30144 18018 0 _0859_
rlabel metal2 29184 18480 29184 18480 0 _0860_
rlabel metal2 29568 18564 29568 18564 0 _0861_
rlabel metal2 32832 19614 32832 19614 0 _0862_
rlabel metal2 32256 19530 32256 19530 0 _0863_
rlabel metal2 32208 18396 32208 18396 0 _0864_
rlabel metal2 32496 19236 32496 19236 0 _0865_
rlabel metal2 36000 19236 36000 19236 0 _0866_
rlabel metal2 35712 19488 35712 19488 0 _0867_
rlabel metal2 35520 19992 35520 19992 0 _0868_
rlabel metal2 35904 20076 35904 20076 0 _0869_
rlabel metal2 37536 19782 37536 19782 0 _0870_
rlabel metal3 38160 19824 38160 19824 0 _0871_
rlabel metal2 38256 19908 38256 19908 0 _0872_
rlabel metal2 38592 21042 38592 21042 0 _0873_
rlabel metal2 43584 18984 43584 18984 0 _0874_
rlabel metal3 42720 18690 42720 18690 0 _0875_
rlabel metal2 41184 20202 41184 20202 0 _0876_
rlabel metal2 42240 19992 42240 19992 0 _0877_
rlabel metal2 44064 16968 44064 16968 0 _0878_
rlabel metal3 42528 17724 42528 17724 0 _0879_
rlabel metal2 42240 18480 42240 18480 0 _0880_
rlabel metal2 41664 17514 41664 17514 0 _0881_
rlabel metal2 42912 13482 42912 13482 0 _0882_
rlabel metal2 42816 13692 42816 13692 0 _0883_
rlabel metal2 41856 14238 41856 14238 0 _0884_
rlabel metal2 41520 13188 41520 13188 0 _0885_
rlabel metal2 39072 15624 39072 15624 0 _0886_
rlabel metal3 39888 15540 39888 15540 0 _0887_
rlabel metal2 40032 14154 40032 14154 0 _0888_
rlabel metal2 39456 14280 39456 14280 0 _0889_
rlabel metal2 36576 16296 36576 16296 0 _0890_
rlabel metal3 37152 16212 37152 16212 0 _0891_
rlabel metal3 38112 14196 38112 14196 0 _0892_
rlabel metal2 36288 15078 36288 15078 0 _0893_
rlabel metal2 34560 16296 34560 16296 0 _0894_
rlabel metal2 34608 16464 34608 16464 0 _0895_
rlabel metal2 34080 15456 34080 15456 0 _0896_
rlabel metal2 33696 15540 33696 15540 0 _0897_
rlabel metal2 32352 13482 32352 13482 0 _0898_
rlabel metal3 32064 13440 32064 13440 0 _0899_
rlabel metal2 32688 13188 32688 13188 0 _0900_
rlabel metal2 32976 13188 32976 13188 0 _0901_
rlabel metal2 36384 13146 36384 13146 0 _0902_
rlabel metal2 36672 11928 36672 11928 0 _0903_
rlabel metal2 35088 12348 35088 12348 0 _0904_
rlabel metal3 35088 11676 35088 11676 0 _0905_
rlabel metal2 38304 11760 38304 11760 0 _0906_
rlabel metal2 38208 11550 38208 11550 0 _0907_
rlabel metal2 36336 11004 36336 11004 0 _0908_
rlabel metal2 36768 11004 36768 11004 0 _0909_
rlabel metal2 42432 10920 42432 10920 0 _0910_
rlabel metal3 41280 10752 41280 10752 0 _0911_
rlabel metal2 39936 9408 39936 9408 0 _0912_
rlabel metal3 40416 9492 40416 9492 0 _0913_
rlabel metal2 44352 10248 44352 10248 0 _0914_
rlabel metal2 42240 9786 42240 9786 0 _0915_
rlabel metal2 42144 9408 42144 9408 0 _0916_
rlabel metal2 42528 9492 42528 9492 0 _0917_
rlabel metal2 46080 9408 46080 9408 0 _0918_
rlabel metal3 45456 9240 45456 9240 0 _0919_
rlabel metal2 44832 7896 44832 7896 0 _0920_
rlabel metal2 45264 7980 45264 7980 0 _0921_
rlabel metal2 48672 8232 48672 8232 0 _0922_
rlabel metal2 48576 8274 48576 8274 0 _0923_
rlabel metal2 47232 7896 47232 7896 0 _0924_
rlabel metal2 47328 6636 47328 6636 0 _0925_
rlabel metal2 48576 6174 48576 6174 0 _0926_
rlabel metal2 48480 5964 48480 5964 0 _0927_
rlabel metal2 47520 5922 47520 5922 0 _0928_
rlabel metal2 47424 4452 47424 4452 0 _0929_
rlabel metal2 52512 3360 52512 3360 0 _0930_
rlabel metal3 51360 3276 51360 3276 0 _0931_
rlabel metal2 49968 3444 49968 3444 0 _0932_
rlabel metal2 50448 3444 50448 3444 0 _0933_
rlabel metal2 54528 6510 54528 6510 0 _0934_
rlabel metal2 54336 6006 54336 6006 0 _0935_
rlabel metal2 52224 5376 52224 5376 0 _0936_
rlabel metal2 52656 5544 52656 5544 0 _0937_
rlabel metal2 53952 9198 53952 9198 0 _0938_
rlabel metal3 54048 7980 54048 7980 0 _0939_
rlabel metal3 53328 7056 53328 7056 0 _0940_
rlabel metal2 52800 7560 52800 7560 0 _0941_
rlabel metal2 53568 10248 53568 10248 0 _0942_
rlabel metal2 53568 10878 53568 10878 0 _0943_
rlabel metal2 53376 8778 53376 8778 0 _0944_
rlabel metal2 52512 9072 52512 9072 0 _0945_
rlabel metal2 51504 11004 51504 11004 0 _0946_
rlabel metal2 51552 10836 51552 10836 0 _0947_
rlabel metal2 51168 8904 51168 8904 0 _0948_
rlabel metal2 50784 11256 50784 11256 0 _0949_
rlabel metal2 48864 12768 48864 12768 0 _0950_
rlabel metal2 49248 12096 49248 12096 0 _0951_
rlabel metal2 48576 11760 48576 11760 0 _0952_
rlabel metal2 48192 12990 48192 12990 0 _0953_
rlabel metal2 47616 14994 47616 14994 0 _0954_
rlabel metal3 47184 14028 47184 14028 0 _0955_
rlabel metal2 46992 13188 46992 13188 0 _0956_
rlabel metal2 46752 11676 46752 11676 0 _0957_
rlabel metal2 46368 15960 46368 15960 0 _0958_
rlabel metal3 46272 15540 46272 15540 0 _0959_
rlabel metal3 45888 14952 45888 14952 0 _0960_
rlabel metal2 45888 15414 45888 15414 0 _0961_
rlabel metal2 48192 18480 48192 18480 0 _0962_
rlabel metal3 48336 18648 48336 18648 0 _0963_
rlabel metal3 46560 17976 46560 17976 0 _0964_
rlabel metal3 47232 18564 47232 18564 0 _0965_
rlabel metal2 51168 16212 51168 16212 0 _0966_
rlabel metal2 49248 16968 49248 16968 0 _0967_
rlabel metal2 49152 17178 49152 17178 0 _0968_
rlabel metal2 49728 16380 49728 16380 0 _0969_
rlabel metal2 52896 14658 52896 14658 0 _0970_
rlabel metal3 52896 14112 52896 14112 0 _0971_
rlabel metal2 51168 14280 51168 14280 0 _0972_
rlabel metal2 51504 14028 51504 14028 0 _0973_
rlabel metal2 56640 14448 56640 14448 0 _0974_
rlabel metal2 56544 13734 56544 13734 0 _0975_
rlabel metal2 54432 13482 54432 13482 0 _0976_
rlabel metal2 54912 13188 54912 13188 0 _0977_
rlabel metal2 58512 13356 58512 13356 0 _0978_
rlabel metal3 57840 13188 57840 13188 0 _0979_
rlabel metal2 56832 13272 56832 13272 0 _0980_
rlabel metal2 56544 12432 56544 12432 0 _0981_
rlabel metal2 59088 10164 59088 10164 0 _0982_
rlabel metal2 59232 10206 59232 10206 0 _0983_
rlabel metal2 57792 10836 57792 10836 0 _0984_
rlabel metal2 58128 10164 58128 10164 0 _0985_
rlabel metal2 59616 8778 59616 8778 0 _0986_
rlabel metal2 59328 8610 59328 8610 0 _0987_
rlabel metal2 58080 9744 58080 9744 0 _0988_
rlabel metal2 57744 8652 57744 8652 0 _0989_
rlabel metal2 60384 6699 60384 6699 0 _0990_
rlabel metal3 59280 6300 59280 6300 0 _0991_
rlabel metal2 58368 6552 58368 6552 0 _0992_
rlabel metal3 58320 6468 58320 6468 0 _0993_
rlabel metal2 61440 5040 61440 5040 0 _0994_
rlabel metal2 61248 6384 61248 6384 0 _0995_
rlabel metal2 59520 5922 59520 5922 0 _0996_
rlabel metal2 59280 4116 59280 4116 0 _0997_
rlabel metal2 56832 3864 56832 3864 0 _0998_
rlabel metal2 57216 4242 57216 4242 0 _0999_
rlabel metal2 57312 4200 57312 4200 0 _1000_
rlabel metal3 56304 4116 56304 4116 0 _1001_
rlabel metal2 57024 2478 57024 2478 0 _1002_
rlabel metal2 56544 2688 56544 2688 0 _1003_
rlabel metal3 56160 1932 56160 1932 0 _1004_
rlabel metal2 55488 1638 55488 1638 0 _1005_
rlabel metal2 60192 2604 60192 2604 0 _1006_
rlabel metal2 59040 2646 59040 2646 0 _1007_
rlabel metal2 57504 1764 57504 1764 0 _1008_
rlabel metal3 59664 924 59664 924 0 _1009_
rlabel metal2 64704 1176 64704 1176 0 _1010_
rlabel metal2 62304 1176 62304 1176 0 _1011_
rlabel metal2 62208 1176 62208 1176 0 _1012_
rlabel metal2 62592 1092 62592 1092 0 _1013_
rlabel metal2 66336 4662 66336 4662 0 _1014_
rlabel metal2 66336 3402 66336 3402 0 _1015_
rlabel via1 64032 2868 64032 2868 0 _1016_
rlabel metal2 64224 3444 64224 3444 0 _1017_
rlabel metal2 66432 6720 66432 6720 0 _1018_
rlabel metal3 66384 5628 66384 5628 0 _1019_
rlabel metal3 65280 5124 65280 5124 0 _1020_
rlabel metal2 65088 5712 65088 5712 0 _1021_
rlabel metal2 65472 7434 65472 7434 0 _1022_
rlabel metal2 65760 7938 65760 7938 0 _1023_
rlabel metal3 64416 7056 64416 7056 0 _1024_
rlabel metal2 63648 8064 63648 8064 0 _1025_
rlabel metal2 64800 10710 64800 10710 0 _1026_
rlabel metal2 64704 10500 64704 10500 0 _1027_
rlabel metal3 19374 36708 19374 36708 0 clk
rlabel metal2 40032 17766 40032 17766 0 clknet_0_clk
rlabel metal3 60000 1092 60000 1092 0 clknet_2_0__leaf_clk
rlabel metal2 31968 15708 31968 15708 0 clknet_2_1__leaf_clk
rlabel metal2 70176 38262 70176 38262 0 clknet_2_2__leaf_clk
rlabel metal2 72720 38220 72720 38220 0 clknet_2_3__leaf_clk
rlabel metal2 2304 15204 2304 15204 0 clknet_leaf_0_clk
rlabel metal2 54432 14994 54432 14994 0 clknet_leaf_10_clk
rlabel metal3 77952 14028 77952 14028 0 clknet_leaf_11_clk
rlabel metal2 74784 9072 74784 9072 0 clknet_leaf_12_clk
rlabel metal2 78192 1092 78192 1092 0 clknet_leaf_13_clk
rlabel metal2 59136 1512 59136 1512 0 clknet_leaf_14_clk
rlabel metal2 55680 8610 55680 8610 0 clknet_leaf_15_clk
rlabel metal2 41568 16842 41568 16842 0 clknet_leaf_16_clk
rlabel metal3 39168 17052 39168 17052 0 clknet_leaf_17_clk
rlabel metal2 2640 5628 2640 5628 0 clknet_leaf_18_clk
rlabel metal2 24096 18480 24096 18480 0 clknet_leaf_1_clk
rlabel metal2 31104 21924 31104 21924 0 clknet_leaf_2_clk
rlabel metal2 43104 27216 43104 27216 0 clknet_leaf_3_clk
rlabel metal2 41376 30786 41376 30786 0 clknet_leaf_4_clk
rlabel metal2 64272 34356 64272 34356 0 clknet_leaf_5_clk
rlabel metal2 65520 35868 65520 35868 0 clknet_leaf_6_clk
rlabel metal2 73104 37968 73104 37968 0 clknet_leaf_7_clk
rlabel metal3 67488 38178 67488 38178 0 clknet_leaf_8_clk
rlabel metal2 42720 19656 42720 19656 0 clknet_leaf_9_clk
rlabel metal2 23136 19362 23136 19362 0 daisychain\[0\]
rlabel metal2 50688 30114 50688 30114 0 daisychain\[100\]
rlabel metal2 51264 28056 51264 28056 0 daisychain\[101\]
rlabel metal2 51744 25578 51744 25578 0 daisychain\[102\]
rlabel metal3 50592 23184 50592 23184 0 daisychain\[103\]
rlabel metal3 47616 22260 47616 22260 0 daisychain\[104\]
rlabel metal2 44736 21798 44736 21798 0 daisychain\[105\]
rlabel metal3 44496 24360 44496 24360 0 daisychain\[106\]
rlabel metal3 45552 25872 45552 25872 0 daisychain\[107\]
rlabel metal3 44256 28308 44256 28308 0 daisychain\[108\]
rlabel metal3 44592 30660 44592 30660 0 daisychain\[109\]
rlabel metal2 36000 15414 36000 15414 0 daisychain\[10\]
rlabel metal3 42240 31164 42240 31164 0 daisychain\[110\]
rlabel metal2 40896 28602 40896 28602 0 daisychain\[111\]
rlabel metal2 39936 26922 39936 26922 0 daisychain\[112\]
rlabel metal2 39936 24192 39936 24192 0 daisychain\[113\]
rlabel metal2 38880 23730 38880 23730 0 daisychain\[114\]
rlabel metal3 36768 24780 36768 24780 0 daisychain\[115\]
rlabel metal2 34272 25746 34272 25746 0 daisychain\[116\]
rlabel metal3 31968 23688 31968 23688 0 daisychain\[117\]
rlabel metal3 30000 22260 30000 22260 0 daisychain\[118\]
rlabel metal3 26400 20076 26400 20076 0 daisychain\[119\]
rlabel metal2 33744 16044 33744 16044 0 daisychain\[11\]
rlabel metal3 4704 2604 4704 2604 0 daisychain\[120\]
rlabel metal3 1824 3360 1824 3360 0 daisychain\[121\]
rlabel metal2 1584 4956 1584 4956 0 daisychain\[122\]
rlabel metal2 1824 7770 1824 7770 0 daisychain\[123\]
rlabel metal2 2016 9114 2016 9114 0 daisychain\[124\]
rlabel metal2 2016 11256 2016 11256 0 daisychain\[125\]
rlabel metal2 2208 12451 2208 12451 0 daisychain\[126\]
rlabel metal2 1632 13944 1632 13944 0 daisychain\[127\]
rlabel metal2 33024 14437 33024 14437 0 daisychain\[12\]
rlabel metal2 36288 12474 36288 12474 0 daisychain\[13\]
rlabel metal2 38784 10710 38784 10710 0 daisychain\[14\]
rlabel metal2 41856 10416 41856 10416 0 daisychain\[15\]
rlabel metal2 43872 9786 43872 9786 0 daisychain\[16\]
rlabel metal3 46224 7980 46224 7980 0 daisychain\[17\]
rlabel metal3 48096 7392 48096 7392 0 daisychain\[18\]
rlabel metal2 48096 4410 48096 4410 0 daisychain\[19\]
rlabel metal2 27024 17724 27024 17724 0 daisychain\[1\]
rlabel metal2 52032 3570 52032 3570 0 daisychain\[20\]
rlabel metal2 53904 6216 53904 6216 0 daisychain\[21\]
rlabel metal2 53520 7980 53520 7980 0 daisychain\[22\]
rlabel metal3 52320 9954 52320 9954 0 daisychain\[23\]
rlabel metal2 50208 11623 50208 11623 0 daisychain\[24\]
rlabel metal2 47760 13188 47760 13188 0 daisychain\[25\]
rlabel metal2 47040 13986 47040 13986 0 daisychain\[26\]
rlabel metal2 45936 17136 45936 17136 0 daisychain\[27\]
rlabel metal2 48672 18858 48672 18858 0 daisychain\[28\]
rlabel via1 50870 15543 50870 15543 0 daisychain\[29\]
rlabel metal2 31872 18816 31872 18816 0 daisychain\[2\]
rlabel metal2 53376 14280 53376 14280 0 daisychain\[30\]
rlabel metal2 56256 14238 56256 14238 0 daisychain\[31\]
rlabel metal3 57792 12684 57792 12684 0 daisychain\[32\]
rlabel metal3 58656 11172 58656 11172 0 daisychain\[33\]
rlabel metal2 58080 8862 58080 8862 0 daisychain\[34\]
rlabel metal2 59232 7014 59232 7014 0 daisychain\[35\]
rlabel metal3 58608 4116 58608 4116 0 daisychain\[36\]
rlabel metal2 55776 2688 55776 2688 0 daisychain\[37\]
rlabel via2 56544 2100 56544 2100 0 daisychain\[38\]
rlabel metal2 61632 2310 61632 2310 0 daisychain\[39\]
rlabel metal2 32928 19866 32928 19866 0 daisychain\[3\]
rlabel metal2 62976 1008 62976 1008 0 daisychain\[40\]
rlabel metal2 65280 3696 65280 3696 0 daisychain\[41\]
rlabel metal2 65376 6132 65376 6132 0 daisychain\[42\]
rlabel metal2 64416 7686 64416 7686 0 daisychain\[43\]
rlabel metal3 64224 9240 64224 9240 0 daisychain\[44\]
rlabel metal2 62784 11413 62784 11413 0 daisychain\[45\]
rlabel metal3 61824 13188 61824 13188 0 daisychain\[46\]
rlabel metal2 64320 14616 64320 14616 0 daisychain\[47\]
rlabel metal2 70080 14322 70080 14322 0 daisychain\[48\]
rlabel metal3 69264 13188 69264 13188 0 daisychain\[49\]
rlabel metal2 37872 20076 37872 20076 0 daisychain\[4\]
rlabel metal3 69120 10164 69120 10164 0 daisychain\[50\]
rlabel metal2 71136 8148 71136 8148 0 daisychain\[51\]
rlabel metal2 71712 5922 71712 5922 0 daisychain\[52\]
rlabel metal2 68400 1932 68400 1932 0 daisychain\[53\]
rlabel metal2 71424 3738 71424 3738 0 daisychain\[54\]
rlabel metal2 73632 2688 73632 2688 0 daisychain\[55\]
rlabel metal2 76560 2604 76560 2604 0 daisychain\[56\]
rlabel metal3 76368 4284 76368 4284 0 daisychain\[57\]
rlabel metal3 74640 6468 74640 6468 0 daisychain\[58\]
rlabel metal2 75936 8568 75936 8568 0 daisychain\[59\]
rlabel metal2 39360 19362 39360 19362 0 daisychain\[5\]
rlabel metal2 75888 10416 75888 10416 0 daisychain\[60\]
rlabel metal2 74928 11928 74928 11928 0 daisychain\[61\]
rlabel metal3 75456 13188 75456 13188 0 daisychain\[62\]
rlabel metal2 74640 13776 74640 13776 0 daisychain\[63\]
rlabel metal2 75744 25116 75744 25116 0 daisychain\[64\]
rlabel metal3 76272 26796 76272 26796 0 daisychain\[65\]
rlabel metal3 75792 29820 75792 29820 0 daisychain\[66\]
rlabel metal2 76032 30912 76032 30912 0 daisychain\[67\]
rlabel metal2 77088 33684 77088 33684 0 daisychain\[68\]
rlabel metal2 76608 34902 76608 34902 0 daisychain\[69\]
rlabel metal3 42528 19278 42528 19278 0 daisychain\[6\]
rlabel metal2 77280 37716 77280 37716 0 daisychain\[70\]
rlabel metal2 72192 36162 72192 36162 0 daisychain\[71\]
rlabel metal2 70464 34902 70464 34902 0 daisychain\[72\]
rlabel metal2 67392 37128 67392 37128 0 daisychain\[73\]
rlabel metal3 66720 35196 66720 35196 0 daisychain\[74\]
rlabel metal2 66048 32550 66048 32550 0 daisychain\[75\]
rlabel metal2 72000 32466 72000 32466 0 daisychain\[76\]
rlabel metal2 70656 30114 70656 30114 0 daisychain\[77\]
rlabel metal2 70560 29106 70560 29106 0 daisychain\[78\]
rlabel metal2 71328 26250 71328 26250 0 daisychain\[79\]
rlabel metal2 41952 17010 41952 17010 0 daisychain\[7\]
rlabel metal2 65664 26376 65664 26376 0 daisychain\[80\]
rlabel metal2 64032 25830 64032 25830 0 daisychain\[81\]
rlabel metal2 64320 28182 64320 28182 0 daisychain\[82\]
rlabel metal2 63264 29946 63264 29946 0 daisychain\[83\]
rlabel metal2 62688 32970 62688 32970 0 daisychain\[84\]
rlabel metal3 61872 35868 61872 35868 0 daisychain\[85\]
rlabel metal2 63552 37002 63552 37002 0 daisychain\[86\]
rlabel metal3 57984 36708 57984 36708 0 daisychain\[87\]
rlabel metal2 56064 35490 56064 35490 0 daisychain\[88\]
rlabel metal3 59568 33264 59568 33264 0 daisychain\[89\]
rlabel metal2 41280 14448 41280 14448 0 daisychain\[8\]
rlabel metal2 60192 30114 60192 30114 0 daisychain\[90\]
rlabel metal2 59712 28056 59712 28056 0 daisychain\[91\]
rlabel metal2 58080 24654 58080 24654 0 daisychain\[92\]
rlabel metal2 55488 27342 55488 27342 0 daisychain\[93\]
rlabel metal3 55200 29316 55200 29316 0 daisychain\[94\]
rlabel metal2 55344 31164 55344 31164 0 daisychain\[95\]
rlabel metal3 54144 33600 54144 33600 0 daisychain\[96\]
rlabel metal3 49008 34356 49008 34356 0 daisychain\[97\]
rlabel metal3 47664 33180 47664 33180 0 daisychain\[98\]
rlabel metal2 50688 32004 50688 32004 0 daisychain\[99\]
rlabel metal2 39168 14238 39168 14238 0 daisychain\[9\]
rlabel metal2 53675 17294 53675 17294 0 digitalen.g\[0\].u.OUTN
rlabel metal2 53565 17378 53565 17378 0 digitalen.g\[0\].u.OUTP
rlabel metal2 79008 16800 79008 16800 0 digitalen.g\[1\].u.OUTN
rlabel metal2 79488 16380 79488 16380 0 digitalen.g\[1\].u.OUTP
rlabel metal2 79565 22828 79565 22828 0 digitalen.g\[2\].u.OUTN
rlabel metal2 79675 22828 79675 22828 0 digitalen.g\[2\].u.OUTP
rlabel metal2 53565 22774 53565 22774 0 digitalen.g\[3\].u.OUTN
rlabel metal2 53675 22732 53675 22732 0 digitalen.g\[3\].u.OUTP
rlabel metal3 99924 21672 99924 21672 0 i_in
rlabel metal3 99924 19992 99924 19992 0 i_out
rlabel metal2 58608 14868 58608 14868 0 net
rlabel metal2 864 37704 864 37704 0 net1
rlabel metal2 864 11802 864 11802 0 net10
rlabel metal2 42624 18606 42624 18606 0 net100
rlabel metal2 42912 18144 42912 18144 0 net101
rlabel metal2 57312 2646 57312 2646 0 net102
rlabel metal2 53472 6048 53472 6048 0 net103
rlabel metal2 53472 14658 53472 14658 0 net104
rlabel metal2 43104 19530 43104 19530 0 net105
rlabel metal2 41088 21672 41088 21672 0 net106
rlabel metal2 45792 22650 45792 22650 0 net107
rlabel metal2 39552 29232 39552 29232 0 net108
rlabel metal2 57696 26502 57696 26502 0 net109
rlabel metal2 864 12390 864 12390 0 net11
rlabel metal3 55344 33264 55344 33264 0 net110
rlabel metal2 54816 32592 54816 32592 0 net111
rlabel metal2 50016 28896 50016 28896 0 net112
rlabel metal2 41760 28476 41760 28476 0 net113
rlabel metal2 64704 2520 64704 2520 0 net114
rlabel metal2 61872 1092 61872 1092 0 net115
rlabel metal2 59568 12516 59568 12516 0 net116
rlabel metal2 70752 9912 70752 9912 0 net117
rlabel metal3 78048 2436 78048 2436 0 net118
rlabel metal3 77472 9492 77472 9492 0 net119
rlabel metal2 864 13314 864 13314 0 net12
rlabel metal2 76512 9534 76512 9534 0 net120
rlabel metal2 74976 13986 74976 13986 0 net121
rlabel metal2 62016 15414 62016 15414 0 net122
rlabel metal3 61056 33684 61056 33684 0 net123
rlabel metal2 66336 34146 66336 34146 0 net124
rlabel metal2 61104 28560 61104 28560 0 net125
rlabel metal2 74496 24696 74496 24696 0 net126
rlabel metal2 71568 33684 71568 33684 0 net127
rlabel metal2 75936 29715 75936 29715 0 net128
rlabel metal2 69312 36792 69312 36792 0 net129
rlabel metal2 1200 14196 1200 14196 0 net13
rlabel metal2 64032 37830 64032 37830 0 net130
rlabel metal2 42816 27006 42816 27006 0 net131
rlabel metal2 22752 18270 22752 18270 0 net132
rlabel metal2 22272 18060 22272 18060 0 net133
rlabel metal2 2592 14826 2592 14826 0 net134
rlabel metal2 22224 18480 22224 18480 0 net135
rlabel metal2 42864 19236 42864 19236 0 net136
rlabel metal2 46944 15036 46944 15036 0 net137
rlabel metal2 53472 9492 53472 9492 0 net138
rlabel metal2 57792 13188 57792 13188 0 net139
rlabel metal2 864 15036 864 15036 0 net14
rlabel metal3 46464 32340 46464 32340 0 net140
rlabel metal3 57264 34356 57264 34356 0 net141
rlabel metal3 55152 33348 55152 33348 0 net142
rlabel metal2 41760 29232 41760 29232 0 net143
rlabel metal2 60384 4326 60384 4326 0 net144
rlabel metal2 61728 13566 61728 13566 0 net145
rlabel metal2 67968 2100 67968 2100 0 net146
rlabel metal2 75456 13104 75456 13104 0 net147
rlabel metal3 66720 34482 66720 34482 0 net148
rlabel metal2 63024 35196 63024 35196 0 net149
rlabel metal2 1248 2730 1248 2730 0 net15
rlabel metal2 71040 35364 71040 35364 0 net150
rlabel metal2 72768 35532 72768 35532 0 net151
rlabel metal2 60768 14742 60768 14742 0 net152
rlabel metal2 21984 19446 21984 19446 0 net153
rlabel metal2 6816 14532 6816 14532 0 net154
rlabel metal2 24192 18228 24192 18228 0 net155
rlabel metal3 24672 18480 24672 18480 0 net156
rlabel metal3 2976 23100 2976 23100 0 net157
rlabel metal2 39264 15456 39264 15456 0 net158
rlabel metal2 42624 12180 42624 12180 0 net159
rlabel metal2 912 2688 912 2688 0 net16
rlabel metal2 56832 2742 56832 2742 0 net160
rlabel metal2 56448 13944 56448 13944 0 net161
rlabel metal3 50496 19992 50496 19992 0 net162
rlabel metal2 37728 22386 37728 22386 0 net163
rlabel metal2 42336 29904 42336 29904 0 net164
rlabel metal2 55008 26082 55008 26082 0 net165
rlabel metal3 52128 35868 52128 35868 0 net166
rlabel metal3 41328 26292 41328 26292 0 net167
rlabel metal2 59808 9324 59808 9324 0 net168
rlabel metal2 62592 14490 62592 14490 0 net169
rlabel metal2 1248 4452 1248 4452 0 net17
rlabel metal2 77472 3318 77472 3318 0 net170
rlabel metal2 76320 11088 76320 11088 0 net171
rlabel metal3 67104 35280 67104 35280 0 net172
rlabel metal2 64128 35322 64128 35322 0 net173
rlabel metal2 72576 35784 72576 35784 0 net174
rlabel metal2 74256 35868 74256 35868 0 net175
rlabel metal4 61920 14910 61920 14910 0 net176
rlabel metal2 1824 23940 1824 23940 0 net177
rlabel metal2 1728 15960 1728 15960 0 net178
rlabel metal2 26496 18354 26496 18354 0 net179
rlabel metal2 816 4200 816 4200 0 net18
rlabel metal2 32496 25284 32496 25284 0 net180
rlabel metal2 22368 20664 22368 20664 0 net181
rlabel metal3 41472 14490 41472 14490 0 net182
rlabel metal2 47520 18480 47520 18480 0 net183
rlabel metal2 55680 4158 55680 4158 0 net184
rlabel metal2 41568 18186 41568 18186 0 net185
rlabel metal2 42336 20328 42336 20328 0 net186
rlabel metal2 42624 30366 42624 30366 0 net187
rlabel metal2 55872 35658 55872 35658 0 net188
rlabel metal2 50688 35028 50688 35028 0 net189
rlabel metal2 912 4872 912 4872 0 net19
rlabel metal2 42432 29652 42432 29652 0 net190
rlabel metal2 60480 1386 60480 1386 0 net191
rlabel metal3 62448 13272 62448 13272 0 net192
rlabel metal2 69696 9786 69696 9786 0 net193
rlabel metal2 74880 13074 74880 13074 0 net194
rlabel metal2 65952 35112 65952 35112 0 net195
rlabel metal2 57312 38094 57312 38094 0 net196
rlabel metal3 68016 37632 68016 37632 0 net197
rlabel metal2 67584 37716 67584 37716 0 net198
rlabel metal2 67824 38052 67824 38052 0 net199
rlabel metal2 864 22218 864 22218 0 net2
rlabel metal2 816 7224 816 7224 0 net20
rlabel metal3 27360 20664 27360 20664 0 net200
rlabel metal2 72672 14700 72672 14700 0 net201
rlabel metal2 68544 24780 68544 24780 0 net202
rlabel metal2 72144 13356 72144 13356 0 net203
rlabel metal2 57552 16380 57552 16380 0 net204
rlabel metal2 72960 11256 72960 11256 0 net205
rlabel metal2 51360 21252 51360 21252 0 net206
rlabel metal2 73920 9744 73920 9744 0 net207
rlabel metal2 53616 16380 53616 16380 0 net208
rlabel metal2 74304 8400 74304 8400 0 net209
rlabel metal2 960 7896 960 7896 0 net21
rlabel metal2 71232 24864 71232 24864 0 net210
rlabel metal3 75216 6300 75216 6300 0 net211
rlabel metal2 50784 18060 50784 18060 0 net212
rlabel metal3 74688 4788 74688 4788 0 net213
rlabel metal2 36192 25956 36192 25956 0 net214
rlabel metal2 76032 2352 76032 2352 0 net215
rlabel metal2 50064 19908 50064 19908 0 net216
rlabel metal2 70944 2352 70944 2352 0 net217
rlabel metal2 71904 27888 71904 27888 0 net218
rlabel metal2 69456 4788 69456 4788 0 net219
rlabel metal3 1152 13776 1152 13776 0 net22
rlabel metal2 46848 16716 46848 16716 0 net220
rlabel metal2 66528 1932 66528 1932 0 net221
rlabel metal2 52608 24108 52608 24108 0 net222
rlabel metal2 69408 6888 69408 6888 0 net223
rlabel metal2 48432 15372 48432 15372 0 net224
rlabel metal2 68544 8358 68544 8358 0 net225
rlabel metal2 72240 31500 72240 31500 0 net226
rlabel metal3 67584 10332 67584 10332 0 net227
rlabel metal2 49824 13074 49824 13074 0 net228
rlabel metal2 67584 12180 67584 12180 0 net229
rlabel metal2 26592 18648 26592 18648 0 net23
rlabel metal2 5520 4788 5520 4788 0 net230
rlabel metal2 68064 15036 68064 15036 0 net231
rlabel metal2 52512 12180 52512 12180 0 net232
rlabel metal2 65136 13356 65136 13356 0 net233
rlabel metal2 72864 32424 72864 32424 0 net234
rlabel metal3 62064 13356 62064 13356 0 net235
rlabel metal2 54336 10668 54336 10668 0 net236
rlabel metal2 62160 11844 62160 11844 0 net237
rlabel metal2 52848 25956 52848 25956 0 net238
rlabel metal2 62400 9912 62400 9912 0 net239
rlabel metal2 32064 24906 32064 24906 0 net24
rlabel metal2 54912 8988 54912 8988 0 net240
rlabel metal2 63024 7812 63024 7812 0 net241
rlabel metal2 67296 31836 67296 31836 0 net242
rlabel metal2 63456 6258 63456 6258 0 net243
rlabel metal2 55104 6888 55104 6888 0 net244
rlabel metal2 63264 3906 63264 3906 0 net245
rlabel metal3 35904 22428 35904 22428 0 net246
rlabel metal2 62208 2352 62208 2352 0 net247
rlabel metal2 52896 4452 52896 4452 0 net248
rlabel metal3 60240 1260 60240 1260 0 net249
rlabel metal2 1728 4872 1728 4872 0 net25
rlabel metal2 67920 34524 67920 34524 0 net250
rlabel metal2 53952 2352 53952 2352 0 net251
rlabel metal2 49344 5796 49344 5796 0 net252
rlabel metal2 55104 4032 55104 4032 0 net253
rlabel metal2 52512 28308 52512 28308 0 net254
rlabel metal2 59712 5376 59712 5376 0 net255
rlabel metal2 49344 7980 49344 7980 0 net256
rlabel metal2 57264 6300 57264 6300 0 net257
rlabel metal2 69696 36960 69696 36960 0 net258
rlabel metal2 56448 8652 56448 8652 0 net259
rlabel via2 41376 16884 41376 16884 0 net26
rlabel metal2 47184 9324 47184 9324 0 net260
rlabel metal2 56352 11634 56352 11634 0 net261
rlabel metal3 5664 12348 5664 12348 0 net262
rlabel metal2 55344 11844 55344 11844 0 net263
rlabel metal3 44736 11844 44736 11844 0 net264
rlabel metal2 54336 14448 54336 14448 0 net265
rlabel metal3 72672 35028 72672 35028 0 net266
rlabel metal2 51024 13860 51024 13860 0 net267
rlabel metal2 42768 12348 42768 12348 0 net268
rlabel metal2 49104 15372 49104 15372 0 net269
rlabel metal2 47616 18648 47616 18648 0 net27
rlabel metal3 51984 30492 51984 30492 0 net270
rlabel metal2 46800 19908 46800 19908 0 net271
rlabel metal2 39552 13158 39552 13158 0 net272
rlabel metal2 43776 15792 43776 15792 0 net273
rlabel metal2 74064 38052 74064 38052 0 net274
rlabel metal2 45120 14448 45120 14448 0 net275
rlabel metal2 37344 13074 37344 13074 0 net276
rlabel metal2 45936 11844 45936 11844 0 net277
rlabel metal3 41760 22932 41760 22932 0 net278
rlabel metal2 48048 10836 48048 10836 0 net279
rlabel metal2 55776 4032 55776 4032 0 net28
rlabel metal2 30432 14280 30432 14280 0 net280
rlabel metal2 50400 9744 50400 9744 0 net281
rlabel metal2 78528 37464 78528 37464 0 net282
rlabel metal2 50976 8379 50976 8379 0 net283
rlabel metal2 34752 17472 34752 17472 0 net284
rlabel metal2 51936 6888 51936 6888 0 net285
rlabel metal2 51600 33012 51600 33012 0 net286
rlabel metal2 50112 4452 50112 4452 0 net287
rlabel metal2 37776 17892 37776 17892 0 net288
rlabel metal2 46176 5376 46176 5376 0 net289
rlabel metal2 41088 17136 41088 17136 0 net29
rlabel metal2 77856 35616 77856 35616 0 net290
rlabel metal2 45888 7476 45888 7476 0 net291
rlabel metal2 40896 15792 40896 15792 0 net292
rlabel metal2 44688 9324 44688 9324 0 net293
rlabel metal2 5856 4788 5856 4788 0 net294
rlabel metal2 41472 8988 41472 8988 0 net295
rlabel metal2 43872 13776 43872 13776 0 net296
rlabel metal2 39840 10500 39840 10500 0 net297
rlabel metal2 77856 33318 77856 33318 0 net298
rlabel metal3 36480 10836 36480 10836 0 net299
rlabel metal2 1488 22932 1488 22932 0 net3
rlabel metal2 42432 19992 42432 19992 0 net30
rlabel metal2 43632 16884 43632 16884 0 net300
rlabel metal2 34320 11844 34320 11844 0 net301
rlabel metal2 46272 33318 46272 33318 0 net302
rlabel metal2 33456 14868 33456 14868 0 net303
rlabel metal3 44448 19908 44448 19908 0 net304
rlabel metal2 31488 15792 31488 15792 0 net305
rlabel metal2 77856 31080 77856 31080 0 net306
rlabel metal3 36288 14868 36288 14868 0 net307
rlabel metal3 39936 19404 39936 19404 0 net308
rlabel metal2 38208 15162 38208 15162 0 net309
rlabel metal2 42528 32088 42528 32088 0 net31
rlabel metal2 41328 25452 41328 25452 0 net310
rlabel metal2 40752 13356 40752 13356 0 net311
rlabel metal2 36672 17892 36672 17892 0 net312
rlabel metal2 40320 19362 40320 19362 0 net313
rlabel metal2 77520 29988 77520 29988 0 net314
rlabel metal2 41808 20916 41808 20916 0 net315
rlabel metal2 33888 18858 33888 18858 0 net316
rlabel metal2 39552 21084 39552 21084 0 net317
rlabel metal2 52512 35196 52512 35196 0 net318
rlabel metal2 35808 21084 35808 21084 0 net319
rlabel metal2 55872 35364 55872 35364 0 net32
rlabel metal2 30816 17502 30816 17502 0 net320
rlabel metal2 32784 21420 32784 21420 0 net321
rlabel metal2 77568 27132 77568 27132 0 net322
rlabel metal2 29712 19908 29712 19908 0 net323
rlabel metal2 27696 17892 27696 17892 0 net324
rlabel metal2 25920 19362 25920 19362 0 net325
rlabel metal2 23280 19908 23280 19908 0 net326
rlabel metal2 23520 17502 23520 17502 0 net327
rlabel metal2 77184 24864 77184 24864 0 net328
rlabel metal2 1488 16380 1488 16380 0 net329
rlabel metal2 53760 32970 53760 32970 0 net33
rlabel metal2 56160 33318 56160 33318 0 net330
rlabel metal2 2496 12768 2496 12768 0 net331
rlabel metal2 76704 15036 76704 15036 0 net332
rlabel metal2 1872 11844 1872 11844 0 net333
rlabel metal2 42240 26376 42240 26376 0 net334
rlabel metal2 1344 8988 1344 8988 0 net335
rlabel metal2 77424 13356 77424 13356 0 net336
rlabel metal2 1632 7476 1632 7476 0 net337
rlabel metal2 56592 32004 56592 32004 0 net338
rlabel metal2 1728 5964 1728 5964 0 net339
rlabel metal4 41184 28644 41184 28644 0 net34
rlabel metal2 77328 11844 77328 11844 0 net340
rlabel metal2 1776 4284 1776 4284 0 net341
rlabel metal2 9792 18816 9792 18816 0 net342
rlabel metal3 7296 19404 7296 19404 0 net343
rlabel metal2 77664 10500 77664 10500 0 net344
rlabel metal2 27840 21084 27840 21084 0 net345
rlabel metal2 56640 29568 56640 29568 0 net346
rlabel metal2 28752 23940 28752 23940 0 net347
rlabel metal2 77616 7812 77616 7812 0 net348
rlabel metal2 30336 25032 30336 25032 0 net349
rlabel metal2 62880 1134 62880 1134 0 net35
rlabel metal2 42528 28644 42528 28644 0 net350
rlabel metal2 32736 25788 32736 25788 0 net351
rlabel metal3 77616 7308 77616 7308 0 net352
rlabel metal2 35520 22986 35520 22986 0 net353
rlabel metal2 55584 25032 55584 25032 0 net354
rlabel metal2 38880 22764 38880 22764 0 net355
rlabel metal3 77664 4788 77664 4788 0 net356
rlabel metal2 37680 25956 37680 25956 0 net357
rlabel metal3 5184 10332 5184 10332 0 net358
rlabel metal2 38256 26964 38256 26964 0 net359
rlabel metal2 57312 10626 57312 10626 0 net36
rlabel metal2 78288 2772 78288 2772 0 net360
rlabel metal2 38928 29988 38928 29988 0 net361
rlabel metal2 60864 24864 60864 24864 0 net362
rlabel metal2 40608 31668 40608 31668 0 net363
rlabel metal3 74304 2772 74304 2772 0 net364
rlabel metal2 44448 30156 44448 30156 0 net365
rlabel metal2 43968 32592 43968 32592 0 net366
rlabel metal2 44736 28476 44736 28476 0 net367
rlabel metal2 72384 4452 72384 4452 0 net368
rlabel metal2 43920 25452 43920 25452 0 net369
rlabel metal2 68352 2562 68352 2562 0 net37
rlabel metal2 61056 26964 61056 26964 0 net370
rlabel metal2 42768 25452 42768 25452 0 net371
rlabel metal2 69408 1596 69408 1596 0 net372
rlabel metal2 42816 22260 42816 22260 0 net373
rlabel metal2 29856 21084 29856 21084 0 net374
rlabel metal2 48144 22428 48144 22428 0 net375
rlabel metal2 72432 7308 72432 7308 0 net376
rlabel metal2 48480 24108 48480 24108 0 net377
rlabel metal2 61104 31500 61104 31500 0 net378
rlabel metal3 48336 25956 48336 25956 0 net379
rlabel metal2 74976 13146 74976 13146 0 net38
rlabel metal2 72144 9324 72144 9324 0 net380
rlabel metal2 49296 28476 49296 28476 0 net381
rlabel metal2 46992 30492 46992 30492 0 net382
rlabel metal2 48384 31080 48384 31080 0 net383
rlabel metal2 71328 10500 71328 10500 0 net384
rlabel metal3 48384 33012 48384 33012 0 net385
rlabel metal2 59184 32844 59184 32844 0 net386
rlabel metal3 46272 34524 46272 34524 0 net387
rlabel metal2 71040 13158 71040 13158 0 net388
rlabel metal3 49824 36036 49824 36036 0 net389
rlabel metal2 66048 35448 66048 35448 0 net39
rlabel metal3 5856 13356 5856 13356 0 net390
rlabel metal2 52752 34524 52752 34524 0 net391
rlabel metal2 71328 15246 71328 15246 0 net392
rlabel metal2 53280 30723 53280 30723 0 net393
rlabel metal3 56256 34524 56256 34524 0 net394
rlabel metal2 53280 29088 53280 29088 0 net395
rlabel metal2 65904 14868 65904 14868 0 net396
rlabel metal2 56208 27468 56208 27468 0 net397
rlabel metal2 47568 28476 47568 28476 0 net398
rlabel metal2 57936 25956 57936 25956 0 net399
rlabel metal3 1440 23856 1440 23856 0 net4
rlabel metal3 62448 32844 62448 32844 0 net40
rlabel metal2 61056 15960 61056 15960 0 net400
rlabel metal2 57744 28476 57744 28476 0 net401
rlabel metal2 60192 37716 60192 37716 0 net402
rlabel metal2 58272 30324 58272 30324 0 net403
rlabel metal2 65280 11844 65280 11844 0 net404
rlabel metal2 58656 34692 58656 34692 0 net405
rlabel metal2 33216 21840 33216 21840 0 net406
rlabel metal2 54912 37128 54912 37128 0 net407
rlabel metal2 65856 10500 65856 10500 0 net408
rlabel metal2 56448 37716 56448 37716 0 net409
rlabel metal2 68160 37830 68160 37830 0 net41
rlabel metal2 64608 37746 64608 37746 0 net410
rlabel metal2 61920 37716 61920 37716 0 net411
rlabel metal2 66480 8820 66480 8820 0 net412
rlabel metal2 60240 36036 60240 36036 0 net413
rlabel metal2 47616 24864 47616 24864 0 net414
rlabel metal3 61056 33012 61056 33012 0 net415
rlabel metal2 67200 6132 67200 6132 0 net416
rlabel metal2 63600 31500 63600 31500 0 net417
rlabel metal2 63552 34692 63552 34692 0 net418
rlabel metal2 62352 28980 62352 28980 0 net419
rlabel metal2 72864 35406 72864 35406 0 net42
rlabel metal2 66864 4788 66864 4788 0 net420
rlabel metal2 62112 26544 62112 26544 0 net421
rlabel metal2 5520 7308 5520 7308 0 net422
rlabel metal2 66432 26376 66432 26376 0 net423
rlabel metal2 65088 1596 65088 1596 0 net424
rlabel metal2 69408 27132 69408 27132 0 net425
rlabel metal2 63696 33516 63696 33516 0 net426
rlabel metal3 67776 28980 67776 28980 0 net427
rlabel metal2 60144 4284 60144 4284 0 net428
rlabel metal3 68736 31500 68736 31500 0 net429
rlabel metal2 74304 15078 74304 15078 0 net43
rlabel metal2 46896 23940 46896 23940 0 net430
rlabel metal2 69744 33516 69744 33516 0 net431
rlabel metal2 57408 1596 57408 1596 0 net432
rlabel metal2 66624 34104 66624 34104 0 net433
rlabel metal2 66480 30492 66480 30492 0 net434
rlabel metal2 64752 35028 64752 35028 0 net435
rlabel metal2 56640 5376 56640 5376 0 net436
rlabel metal2 66240 37746 66240 37746 0 net437
rlabel metal2 33600 22986 33600 22986 0 net438
rlabel metal2 69504 36078 69504 36078 0 net439
rlabel metal2 2208 16002 2208 16002 0 net44
rlabel metal2 61728 5964 61728 5964 0 net440
rlabel metal3 72480 37044 72480 37044 0 net441
rlabel metal2 66240 27888 66240 27888 0 net442
rlabel metal2 75984 38052 75984 38052 0 net443
rlabel metal2 60960 8400 60960 8400 0 net444
rlabel metal2 74640 36036 74640 36036 0 net445
rlabel metal2 46464 22008 46464 22008 0 net446
rlabel metal2 75024 33516 75024 33516 0 net447
rlabel metal2 60288 10164 60288 10164 0 net448
rlabel metal2 74064 32004 74064 32004 0 net449
rlabel metal2 25632 19194 25632 19194 0 net45
rlabel metal2 64800 24864 64800 24864 0 net450
rlabel metal2 73920 29568 73920 29568 0 net451
rlabel metal2 59760 12348 59760 12348 0 net452
rlabel metal2 73536 27300 73536 27300 0 net453
rlabel metal2 5040 15372 5040 15372 0 net454
rlabel metal2 73536 25452 73536 25452 0 net455
rlabel metal3 366 15708 366 15708 0 net456
rlabel metal3 366 16548 366 16548 0 net457
rlabel metal3 366 17388 366 17388 0 net458
rlabel metal3 366 18228 366 18228 0 net459
rlabel metal2 26688 20538 26688 20538 0 net46
rlabel metal3 366 19068 366 19068 0 net460
rlabel metal3 366 19908 366 19908 0 net461
rlabel metal3 366 20748 366 20748 0 net462
rlabel metal3 366 21588 366 21588 0 net463
rlabel metal3 26544 19992 26544 19992 0 net47
rlabel metal3 2736 2604 2736 2604 0 net48
rlabel metal2 40128 13944 40128 13944 0 net49
rlabel metal3 1824 25116 1824 25116 0 net5
rlabel metal2 56064 2541 56064 2541 0 net50
rlabel metal2 53664 14826 53664 14826 0 net51
rlabel metal2 41952 19068 41952 19068 0 net52
rlabel metal2 41808 22932 41808 22932 0 net53
rlabel metal3 57600 35196 57600 35196 0 net54
rlabel metal2 54144 33138 54144 33138 0 net55
rlabel metal2 41664 29946 41664 29946 0 net56
rlabel metal2 62016 1050 62016 1050 0 net57
rlabel metal2 58752 10290 58752 10290 0 net58
rlabel metal2 76176 2604 76176 2604 0 net59
rlabel metal3 4032 25956 4032 25956 0 net6
rlabel metal2 75648 8484 75648 8484 0 net60
rlabel metal2 66144 33978 66144 33978 0 net61
rlabel metal2 67104 36792 67104 36792 0 net62
rlabel metal2 71904 35994 71904 35994 0 net63
rlabel metal2 60048 36708 60048 36708 0 net64
rlabel metal2 74784 14406 74784 14406 0 net65
rlabel metal2 25920 21294 25920 21294 0 net66
rlabel metal3 22176 17724 22176 17724 0 net67
rlabel metal2 33600 16548 33600 16548 0 net68
rlabel metal2 21888 18270 21888 18270 0 net69
rlabel metal2 1536 17418 1536 17418 0 net7
rlabel metal2 6336 4872 6336 4872 0 net70
rlabel metal3 42432 14700 42432 14700 0 net71
rlabel metal3 47088 16800 47088 16800 0 net72
rlabel metal2 55680 4872 55680 4872 0 net73
rlabel metal2 56928 14616 56928 14616 0 net74
rlabel metal2 46560 31374 46560 31374 0 net75
rlabel metal3 58656 34608 58656 34608 0 net76
rlabel metal2 55488 32130 55488 32130 0 net77
rlabel metal3 41424 22848 41424 22848 0 net78
rlabel metal2 58896 2604 58896 2604 0 net79
rlabel metal3 1200 9660 1200 9660 0 net8
rlabel metal2 60960 14490 60960 14490 0 net80
rlabel metal3 77616 2184 77616 2184 0 net81
rlabel metal2 76992 7896 76992 7896 0 net82
rlabel metal2 60192 25788 60192 25788 0 net83
rlabel metal2 63600 38220 63600 38220 0 net84
rlabel metal2 69168 37548 69168 37548 0 net85
rlabel metal2 76224 25116 76224 25116 0 net86
rlabel metal3 61632 14868 61632 14868 0 net87
rlabel metal2 22080 20748 22080 20748 0 net88
rlabel metal2 3264 2730 3264 2730 0 net89
rlabel metal2 864 10878 864 10878 0 net9
rlabel metal2 4800 8736 4800 8736 0 net90
rlabel metal2 31968 19572 31968 19572 0 net91
rlabel metal2 38496 13986 38496 13986 0 net92
rlabel metal2 25440 18312 25440 18312 0 net93
rlabel metal2 32256 20790 32256 20790 0 net94
rlabel metal2 36528 22596 36528 22596 0 net95
rlabel metal2 26880 19992 26880 19992 0 net96
rlabel metal2 24384 18438 24384 18438 0 net97
rlabel metal2 42336 9954 42336 9954 0 net98
rlabel metal2 49536 12390 49536 12390 0 net99
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal2 25536 17598 25536 17598 0 state\[0\]
rlabel metal2 54336 27090 54336 27090 0 state\[100\]
rlabel metal2 54720 26502 54720 26502 0 state\[101\]
rlabel metal2 54816 25032 54816 25032 0 state\[102\]
rlabel metal2 54144 23646 54144 23646 0 state\[103\]
rlabel metal2 63275 22828 63275 22828 0 state\[104\]
rlabel metal2 62875 22828 62875 22828 0 state\[105\]
rlabel metal2 62475 22828 62475 22828 0 state\[106\]
rlabel metal2 62075 22828 62075 22828 0 state\[107\]
rlabel metal2 61675 22828 61675 22828 0 state\[108\]
rlabel metal2 61275 22828 61275 22828 0 state\[109\]
rlabel metal4 39744 16758 39744 16758 0 state\[10\]
rlabel metal2 43104 31080 43104 31080 0 state\[110\]
rlabel metal2 44352 27972 44352 27972 0 state\[111\]
rlabel metal2 41568 26712 41568 26712 0 state\[112\]
rlabel metal2 41088 24570 41088 24570 0 state\[113\]
rlabel metal3 41424 21672 41424 21672 0 state\[114\]
rlabel metal3 40656 22428 40656 22428 0 state\[115\]
rlabel metal2 38112 26502 38112 26502 0 state\[116\]
rlabel metal3 32736 23772 32736 23772 0 state\[117\]
rlabel metal2 32064 21714 32064 21714 0 state\[118\]
rlabel metal3 32064 21000 32064 21000 0 state\[119\]
rlabel metal2 34368 17304 34368 17304 0 state\[11\]
rlabel metal2 56875 22828 56875 22828 0 state\[120\]
rlabel metal3 56317 23016 56317 23016 0 state\[121\]
rlabel metal2 56069 22764 56069 22764 0 state\[122\]
rlabel metal2 55675 22828 55675 22828 0 state\[123\]
rlabel metal2 55275 22690 55275 22690 0 state\[124\]
rlabel metal2 1440 13146 1440 13146 0 state\[125\]
rlabel metal3 54453 22764 54453 22764 0 state\[126\]
rlabel metal2 36192 16632 36192 16632 0 state\[127\]
rlabel metal2 32448 14280 32448 14280 0 state\[12\]
rlabel metal2 39360 13062 39360 13062 0 state\[13\]
rlabel metal2 59565 17294 59565 17294 0 state\[14\]
rlabel metal2 59965 17294 59965 17294 0 state\[15\]
rlabel metal2 60365 17252 60365 17252 0 state\[16\]
rlabel metal2 60480 16212 60480 16212 0 state\[17\]
rlabel metal2 61440 16128 61440 16128 0 state\[18\]
rlabel metal2 62112 16044 62112 16044 0 state\[19\]
rlabel metal2 27168 17514 27168 17514 0 state\[1\]
rlabel metal3 61296 16212 61296 16212 0 state\[20\]
rlabel metal2 62688 16170 62688 16170 0 state\[21\]
rlabel metal2 62976 15876 62976 15876 0 state\[22\]
rlabel metal2 63264 15834 63264 15834 0 state\[23\]
rlabel metal3 56064 15960 56064 15960 0 state\[24\]
rlabel metal3 57504 13398 57504 13398 0 state\[25\]
rlabel metal2 50400 15162 50400 15162 0 state\[26\]
rlabel metal3 51456 16926 51456 16926 0 state\[27\]
rlabel metal2 52032 18774 52032 18774 0 state\[28\]
rlabel metal2 53856 16884 53856 16884 0 state\[29\]
rlabel metal2 32832 17430 32832 17430 0 state\[2\]
rlabel metal3 59424 15456 59424 15456 0 state\[30\]
rlabel metal2 59520 15834 59520 15834 0 state\[31\]
rlabel metal2 60624 13776 60624 13776 0 state\[32\]
rlabel metal2 61728 12264 61728 12264 0 state\[33\]
rlabel metal2 60192 8946 60192 8946 0 state\[34\]
rlabel metal2 60096 8064 60096 8064 0 state\[35\]
rlabel metal2 62016 5334 62016 5334 0 state\[36\]
rlabel metal2 56448 4410 56448 4410 0 state\[37\]
rlabel metal2 59040 1554 59040 1554 0 state\[38\]
rlabel metal2 59616 2604 59616 2604 0 state\[39\]
rlabel metal2 33504 17976 33504 17976 0 state\[3\]
rlabel metal2 65040 2604 65040 2604 0 state\[40\]
rlabel metal2 70365 17336 70365 17336 0 state\[41\]
rlabel metal2 70765 17294 70765 17294 0 state\[42\]
rlabel metal2 70944 15918 70944 15918 0 state\[43\]
rlabel metal2 71424 16212 71424 16212 0 state\[44\]
rlabel metal2 71965 17294 71965 17294 0 state\[45\]
rlabel metal2 62400 14406 62400 14406 0 state\[46\]
rlabel metal2 72576 16674 72576 16674 0 state\[47\]
rlabel metal2 72960 16674 72960 16674 0 state\[48\]
rlabel metal2 73565 17336 73565 17336 0 state\[49\]
rlabel metal2 38592 18102 38592 18102 0 state\[4\]
rlabel metal2 73632 16212 73632 16212 0 state\[50\]
rlabel metal2 74352 16212 74352 16212 0 state\[51\]
rlabel metal2 74592 15078 74592 15078 0 state\[52\]
rlabel metal2 74976 16674 74976 16674 0 state\[53\]
rlabel metal3 75120 16212 75120 16212 0 state\[54\]
rlabel metal3 74544 2604 74544 2604 0 state\[55\]
rlabel metal2 77088 1974 77088 1974 0 state\[56\]
rlabel metal2 76992 16002 76992 16002 0 state\[57\]
rlabel metal3 77424 16212 77424 16212 0 state\[58\]
rlabel metal2 77424 16212 77424 16212 0 state\[59\]
rlabel metal2 41184 18690 41184 18690 0 state\[5\]
rlabel metal2 77904 16212 77904 16212 0 state\[60\]
rlabel metal2 78288 16212 78288 16212 0 state\[61\]
rlabel metal2 78624 16674 78624 16674 0 state\[62\]
rlabel metal2 79200 16632 79200 16632 0 state\[63\]
rlabel metal2 79275 22828 79275 22828 0 state\[64\]
rlabel metal3 78749 22764 78749 22764 0 state\[65\]
rlabel metal2 78453 22848 78453 22848 0 state\[66\]
rlabel metal2 78075 22828 78075 22828 0 state\[67\]
rlabel metal2 77675 22828 77675 22828 0 state\[68\]
rlabel metal3 78816 34356 78816 34356 0 state\[69\]
rlabel metal2 56160 16128 56160 16128 0 state\[6\]
rlabel metal2 76875 22690 76875 22690 0 state\[70\]
rlabel metal2 73056 35910 73056 35910 0 state\[71\]
rlabel metal2 71808 33936 71808 33936 0 state\[72\]
rlabel metal3 71328 37212 71328 37212 0 state\[73\]
rlabel metal2 66720 34902 66720 34902 0 state\[74\]
rlabel metal2 74875 22732 74875 22732 0 state\[75\]
rlabel metal2 74475 22828 74475 22828 0 state\[76\]
rlabel metal2 74075 22828 74075 22828 0 state\[77\]
rlabel metal2 73675 22828 73675 22828 0 state\[78\]
rlabel metal2 73275 22828 73275 22828 0 state\[79\]
rlabel metal3 42720 16212 42720 16212 0 state\[7\]
rlabel metal2 72875 22828 72875 22828 0 state\[80\]
rlabel metal2 72475 22828 72475 22828 0 state\[81\]
rlabel metal2 68160 28098 68160 28098 0 state\[82\]
rlabel metal2 71675 22828 71675 22828 0 state\[83\]
rlabel metal2 71275 22828 71275 22828 0 state\[84\]
rlabel metal2 65472 34146 65472 34146 0 state\[85\]
rlabel metal2 66720 36582 66720 36582 0 state\[86\]
rlabel metal2 69216 36750 69216 36750 0 state\[87\]
rlabel metal2 57984 34902 57984 34902 0 state\[88\]
rlabel metal2 61152 32256 61152 32256 0 state\[89\]
rlabel metal2 56880 16212 56880 16212 0 state\[8\]
rlabel metal2 63072 29442 63072 29442 0 state\[90\]
rlabel metal2 62976 26964 62976 26964 0 state\[91\]
rlabel metal2 60096 24696 60096 24696 0 state\[92\]
rlabel metal2 55968 24906 55968 24906 0 state\[93\]
rlabel metal2 58560 28770 58560 28770 0 state\[94\]
rlabel metal2 58560 31122 58560 31122 0 state\[95\]
rlabel metal2 55104 33684 55104 33684 0 state\[96\]
rlabel metal2 54432 35658 54432 35658 0 state\[97\]
rlabel metal2 48288 32382 48288 32382 0 state\[98\]
rlabel metal2 51264 32760 51264 32760 0 state\[99\]
rlabel metal2 42720 16548 42720 16548 0 state\[9\]
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 25788 366 25788 0 ui_in[4]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 558 14028 558 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 558 2268 558 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 558 3948 558 3948 0 uo_out[2]
rlabel metal2 672 4536 672 4536 0 uo_out[3]
rlabel metal2 672 5376 672 5376 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
