* Extracted by KLayout with SG13G2 LVS runset on : 19/08/2025 02:06

.SUBCKT PCASCSRCREFL
M$1 \$1 \$2 \$5 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$2 \$5 \$3 \$2 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
.ENDS PCASCSRCREFL
