module heichips25_template (analog_pin0,
    analog_pin1,
    analog_pin2,
    analog_pin3,
    clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 inout analog_pin0;
 inout analog_pin1;
 inout analog_pin2;
 inout analog_pin3;
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net;

 sg13g2_tielo heichips25_template_1 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net1));
 sg13g2_tielo heichips25_template_2 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net2));
 sg13g2_tielo heichips25_template_3 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net3));
 sg13g2_tielo heichips25_template_4 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net4));
 sg13g2_tielo heichips25_template_5 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net5));
 sg13g2_tielo heichips25_template_6 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net6));
 sg13g2_tielo heichips25_template_7 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net7));
 sg13g2_tielo heichips25_template_8 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net8));
 sg13g2_tielo heichips25_template_9 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net9));
 sg13g2_tielo heichips25_template_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_tielo heichips25_template_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_template_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_template_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_template_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_template_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_template_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tielo heichips25_template_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_tielo heichips25_template_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo heichips25_template_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo heichips25_template_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo heichips25_template_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo heichips25_template_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tielo heichips25_template_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1022 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net;
 assign uio_out[3] = net1;
 assign uio_out[4] = net2;
 assign uio_out[5] = net3;
 assign uio_out[6] = net4;
 assign uio_out[7] = net5;
 assign uo_out[0] = net6;
 assign uo_out[1] = net7;
 assign uo_out[2] = net8;
 assign uo_out[3] = net9;
 assign uo_out[4] = net10;
 assign uo_out[5] = net11;
 assign uo_out[6] = net12;
 assign uo_out[7] = net13;
endmodule
