module heichips25_template (analog_pin0,
    analog_pin1,
    analog_pin2,
    analog_pin3,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 inout analog_pin0;
 inout analog_pin1;
 inout analog_pin2;
 inout analog_pin3;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net;

 sg13g2_tielo heichips25_template_1 (.L_LO(net1));
 sg13g2_tielo heichips25_template_2 (.L_LO(net2));
 sg13g2_tielo heichips25_template_3 (.L_LO(net3));
 sg13g2_tielo heichips25_template_4 (.L_LO(net4));
 sg13g2_tielo heichips25_template_5 (.L_LO(net5));
 sg13g2_tielo heichips25_template_6 (.L_LO(net6));
 sg13g2_tielo heichips25_template_7 (.L_LO(net7));
 sg13g2_tielo heichips25_template_8 (.L_LO(net8));
 sg13g2_tielo heichips25_template_9 (.L_LO(net9));
 sg13g2_tielo heichips25_template_10 (.L_LO(net10));
 sg13g2_tielo heichips25_template_11 (.L_LO(net11));
 sg13g2_tielo heichips25_template_12 (.L_LO(net12));
 sg13g2_tielo heichips25_template_13 (.L_LO(net13));
 sg13g2_tielo heichips25_template_14 (.L_LO(net14));
 sg13g2_tielo heichips25_template_15 (.L_LO(net15));
 sg13g2_tielo heichips25_template_16 (.L_LO(net16));
 sg13g2_tielo heichips25_template_17 (.L_LO(net17));
 sg13g2_tielo heichips25_template_18 (.L_LO(net18));
 sg13g2_tielo heichips25_template_19 (.L_LO(net19));
 sg13g2_tielo heichips25_template_20 (.L_LO(net20));
 sg13g2_tielo heichips25_template_21 (.L_LO(net21));
 sg13g2_tielo heichips25_template_22 (.L_LO(net22));
 sg13g2_tielo heichips25_template_23 (.L_LO(net23));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo heichips25_template (.L_LO(net));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_564 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_872 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_8 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_942 ();
 sg13g2_decap_8 FILLER_3_949 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_decap_8 FILLER_4_473 ();
 sg13g2_decap_8 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_8 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_501 ();
 sg13g2_decap_8 FILLER_4_508 ();
 sg13g2_decap_8 FILLER_4_515 ();
 sg13g2_decap_8 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_4_529 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_557 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_571 ();
 sg13g2_decap_8 FILLER_4_578 ();
 sg13g2_decap_8 FILLER_4_585 ();
 sg13g2_decap_8 FILLER_4_592 ();
 sg13g2_decap_8 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_620 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_669 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_711 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_8 FILLER_4_732 ();
 sg13g2_decap_8 FILLER_4_739 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_774 ();
 sg13g2_decap_8 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_8 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_8 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_928 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1026 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_decap_8 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_6_865 ();
 sg13g2_decap_8 FILLER_6_872 ();
 sg13g2_decap_8 FILLER_6_879 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_decap_8 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_487 ();
 sg13g2_decap_8 FILLER_8_494 ();
 sg13g2_decap_8 FILLER_8_501 ();
 sg13g2_decap_8 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_decap_8 FILLER_8_543 ();
 sg13g2_decap_8 FILLER_8_550 ();
 sg13g2_decap_8 FILLER_8_557 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_613 ();
 sg13g2_decap_8 FILLER_8_620 ();
 sg13g2_decap_8 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_decap_8 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_decap_8 FILLER_8_879 ();
 sg13g2_decap_8 FILLER_8_886 ();
 sg13g2_decap_8 FILLER_8_893 ();
 sg13g2_decap_8 FILLER_8_900 ();
 sg13g2_decap_8 FILLER_8_907 ();
 sg13g2_decap_8 FILLER_8_914 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_8_928 ();
 sg13g2_decap_8 FILLER_8_935 ();
 sg13g2_decap_8 FILLER_8_942 ();
 sg13g2_decap_8 FILLER_8_949 ();
 sg13g2_decap_8 FILLER_8_956 ();
 sg13g2_decap_8 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_970 ();
 sg13g2_decap_8 FILLER_8_977 ();
 sg13g2_decap_8 FILLER_8_984 ();
 sg13g2_decap_8 FILLER_8_991 ();
 sg13g2_decap_8 FILLER_8_998 ();
 sg13g2_decap_8 FILLER_8_1005 ();
 sg13g2_decap_8 FILLER_8_1012 ();
 sg13g2_decap_8 FILLER_8_1019 ();
 sg13g2_fill_2 FILLER_8_1026 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_564 ();
 sg13g2_decap_8 FILLER_9_571 ();
 sg13g2_decap_8 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_decap_8 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_8 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_872 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_8 FILLER_9_921 ();
 sg13g2_decap_8 FILLER_9_928 ();
 sg13g2_decap_8 FILLER_9_935 ();
 sg13g2_decap_8 FILLER_9_942 ();
 sg13g2_decap_8 FILLER_9_949 ();
 sg13g2_decap_8 FILLER_9_956 ();
 sg13g2_decap_8 FILLER_9_963 ();
 sg13g2_decap_8 FILLER_9_970 ();
 sg13g2_decap_8 FILLER_9_977 ();
 sg13g2_decap_8 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_decap_8 FILLER_9_998 ();
 sg13g2_decap_8 FILLER_9_1005 ();
 sg13g2_decap_8 FILLER_9_1012 ();
 sg13g2_decap_8 FILLER_9_1019 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_564 ();
 sg13g2_decap_8 FILLER_12_571 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_8 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_8 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_8 FILLER_12_935 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_8 FILLER_13_473 ();
 sg13g2_decap_8 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_decap_8 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_543 ();
 sg13g2_decap_8 FILLER_13_550 ();
 sg13g2_decap_8 FILLER_13_557 ();
 sg13g2_decap_8 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_571 ();
 sg13g2_decap_8 FILLER_13_578 ();
 sg13g2_decap_8 FILLER_13_585 ();
 sg13g2_decap_8 FILLER_13_592 ();
 sg13g2_decap_8 FILLER_13_599 ();
 sg13g2_decap_8 FILLER_13_606 ();
 sg13g2_decap_8 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_879 ();
 sg13g2_decap_8 FILLER_13_886 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_914 ();
 sg13g2_decap_8 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_decap_8 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_942 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_decap_8 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_decap_8 FILLER_14_452 ();
 sg13g2_decap_8 FILLER_14_459 ();
 sg13g2_decap_8 FILLER_14_466 ();
 sg13g2_decap_8 FILLER_14_473 ();
 sg13g2_decap_8 FILLER_14_480 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_decap_8 FILLER_14_515 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_decap_8 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_550 ();
 sg13g2_decap_8 FILLER_14_557 ();
 sg13g2_decap_8 FILLER_14_564 ();
 sg13g2_decap_8 FILLER_14_571 ();
 sg13g2_decap_8 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_585 ();
 sg13g2_decap_8 FILLER_14_592 ();
 sg13g2_decap_8 FILLER_14_599 ();
 sg13g2_decap_8 FILLER_14_606 ();
 sg13g2_decap_8 FILLER_14_613 ();
 sg13g2_decap_8 FILLER_14_620 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_634 ();
 sg13g2_decap_8 FILLER_14_641 ();
 sg13g2_decap_8 FILLER_14_648 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_683 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_704 ();
 sg13g2_decap_8 FILLER_14_711 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_774 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_788 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_816 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_8 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_14_865 ();
 sg13g2_decap_8 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_decap_8 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_decap_8 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_942 ();
 sg13g2_decap_8 FILLER_14_949 ();
 sg13g2_decap_8 FILLER_14_956 ();
 sg13g2_decap_8 FILLER_14_963 ();
 sg13g2_decap_8 FILLER_14_970 ();
 sg13g2_decap_8 FILLER_14_977 ();
 sg13g2_decap_8 FILLER_14_984 ();
 sg13g2_decap_8 FILLER_14_991 ();
 sg13g2_decap_8 FILLER_14_998 ();
 sg13g2_decap_8 FILLER_14_1005 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_fill_2 FILLER_14_1026 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_893 ();
 sg13g2_decap_8 FILLER_15_900 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_914 ();
 sg13g2_decap_8 FILLER_15_921 ();
 sg13g2_decap_8 FILLER_15_928 ();
 sg13g2_decap_8 FILLER_15_935 ();
 sg13g2_decap_8 FILLER_15_942 ();
 sg13g2_decap_8 FILLER_15_949 ();
 sg13g2_decap_8 FILLER_15_956 ();
 sg13g2_decap_8 FILLER_15_963 ();
 sg13g2_decap_8 FILLER_15_970 ();
 sg13g2_decap_8 FILLER_15_977 ();
 sg13g2_decap_8 FILLER_15_984 ();
 sg13g2_decap_8 FILLER_15_991 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_decap_8 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_decap_8 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_15_1026 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_decap_8 FILLER_16_438 ();
 sg13g2_decap_8 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_452 ();
 sg13g2_decap_8 FILLER_16_459 ();
 sg13g2_decap_8 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_473 ();
 sg13g2_decap_8 FILLER_16_480 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_decap_8 FILLER_16_494 ();
 sg13g2_decap_8 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_8 FILLER_16_515 ();
 sg13g2_decap_8 FILLER_16_522 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_8 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_613 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_8 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_865 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_decap_8 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_963 ();
 sg13g2_decap_8 FILLER_16_970 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_decap_8 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_991 ();
 sg13g2_decap_8 FILLER_16_998 ();
 sg13g2_decap_8 FILLER_16_1005 ();
 sg13g2_decap_8 FILLER_16_1012 ();
 sg13g2_decap_8 FILLER_16_1019 ();
 sg13g2_fill_2 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_decap_8 FILLER_18_466 ();
 sg13g2_decap_8 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_480 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_543 ();
 sg13g2_decap_8 FILLER_18_550 ();
 sg13g2_decap_8 FILLER_18_557 ();
 sg13g2_decap_8 FILLER_18_564 ();
 sg13g2_decap_8 FILLER_18_571 ();
 sg13g2_decap_8 FILLER_18_578 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_decap_8 FILLER_18_592 ();
 sg13g2_decap_8 FILLER_18_599 ();
 sg13g2_decap_8 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_613 ();
 sg13g2_decap_8 FILLER_18_620 ();
 sg13g2_decap_8 FILLER_18_627 ();
 sg13g2_decap_8 FILLER_18_634 ();
 sg13g2_decap_8 FILLER_18_641 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_655 ();
 sg13g2_decap_8 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_669 ();
 sg13g2_decap_8 FILLER_18_676 ();
 sg13g2_decap_8 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_844 ();
 sg13g2_decap_8 FILLER_18_851 ();
 sg13g2_decap_8 FILLER_18_858 ();
 sg13g2_decap_8 FILLER_18_865 ();
 sg13g2_decap_8 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_879 ();
 sg13g2_decap_8 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_893 ();
 sg13g2_decap_8 FILLER_18_900 ();
 sg13g2_decap_8 FILLER_18_907 ();
 sg13g2_decap_8 FILLER_18_914 ();
 sg13g2_decap_8 FILLER_18_921 ();
 sg13g2_decap_8 FILLER_18_928 ();
 sg13g2_decap_8 FILLER_18_935 ();
 sg13g2_decap_8 FILLER_18_942 ();
 sg13g2_decap_8 FILLER_18_949 ();
 sg13g2_decap_8 FILLER_18_956 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_decap_8 FILLER_18_970 ();
 sg13g2_decap_8 FILLER_18_977 ();
 sg13g2_decap_8 FILLER_18_984 ();
 sg13g2_decap_8 FILLER_18_991 ();
 sg13g2_decap_8 FILLER_18_998 ();
 sg13g2_decap_8 FILLER_18_1005 ();
 sg13g2_decap_8 FILLER_18_1012 ();
 sg13g2_decap_8 FILLER_18_1019 ();
 sg13g2_fill_2 FILLER_18_1026 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_8 FILLER_19_424 ();
 sg13g2_decap_8 FILLER_19_431 ();
 sg13g2_decap_8 FILLER_19_438 ();
 sg13g2_decap_8 FILLER_19_445 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_decap_8 FILLER_19_473 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_decap_8 FILLER_19_487 ();
 sg13g2_decap_8 FILLER_19_494 ();
 sg13g2_decap_8 FILLER_19_501 ();
 sg13g2_decap_8 FILLER_19_508 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_8 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_8 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_19_865 ();
 sg13g2_decap_8 FILLER_19_872 ();
 sg13g2_decap_8 FILLER_19_879 ();
 sg13g2_decap_8 FILLER_19_886 ();
 sg13g2_decap_8 FILLER_19_893 ();
 sg13g2_decap_8 FILLER_19_900 ();
 sg13g2_decap_8 FILLER_19_907 ();
 sg13g2_decap_8 FILLER_19_914 ();
 sg13g2_decap_8 FILLER_19_921 ();
 sg13g2_decap_8 FILLER_19_928 ();
 sg13g2_decap_8 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_942 ();
 sg13g2_decap_8 FILLER_19_949 ();
 sg13g2_decap_8 FILLER_19_956 ();
 sg13g2_decap_8 FILLER_19_963 ();
 sg13g2_decap_8 FILLER_19_970 ();
 sg13g2_decap_8 FILLER_19_977 ();
 sg13g2_decap_8 FILLER_19_984 ();
 sg13g2_decap_8 FILLER_19_991 ();
 sg13g2_decap_8 FILLER_19_998 ();
 sg13g2_decap_8 FILLER_19_1005 ();
 sg13g2_decap_8 FILLER_19_1012 ();
 sg13g2_decap_8 FILLER_19_1019 ();
 sg13g2_fill_2 FILLER_19_1026 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_decap_8 FILLER_20_438 ();
 sg13g2_decap_8 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_466 ();
 sg13g2_decap_8 FILLER_20_473 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_decap_8 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_522 ();
 sg13g2_decap_8 FILLER_20_529 ();
 sg13g2_decap_8 FILLER_20_536 ();
 sg13g2_decap_8 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_decap_8 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_592 ();
 sg13g2_decap_8 FILLER_20_599 ();
 sg13g2_decap_8 FILLER_20_606 ();
 sg13g2_decap_8 FILLER_20_613 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_648 ();
 sg13g2_decap_8 FILLER_20_655 ();
 sg13g2_decap_8 FILLER_20_662 ();
 sg13g2_decap_8 FILLER_20_669 ();
 sg13g2_decap_8 FILLER_20_676 ();
 sg13g2_decap_8 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_decap_8 FILLER_20_697 ();
 sg13g2_decap_8 FILLER_20_704 ();
 sg13g2_decap_8 FILLER_20_711 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_725 ();
 sg13g2_decap_8 FILLER_20_732 ();
 sg13g2_decap_8 FILLER_20_739 ();
 sg13g2_decap_8 FILLER_20_746 ();
 sg13g2_decap_8 FILLER_20_753 ();
 sg13g2_decap_8 FILLER_20_760 ();
 sg13g2_decap_8 FILLER_20_767 ();
 sg13g2_decap_8 FILLER_20_774 ();
 sg13g2_decap_8 FILLER_20_781 ();
 sg13g2_decap_8 FILLER_20_788 ();
 sg13g2_decap_8 FILLER_20_795 ();
 sg13g2_decap_8 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_809 ();
 sg13g2_decap_8 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_8 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_879 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_914 ();
 sg13g2_decap_8 FILLER_20_921 ();
 sg13g2_decap_8 FILLER_20_928 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_decap_8 FILLER_20_942 ();
 sg13g2_decap_8 FILLER_20_949 ();
 sg13g2_decap_8 FILLER_20_956 ();
 sg13g2_decap_8 FILLER_20_963 ();
 sg13g2_decap_8 FILLER_20_970 ();
 sg13g2_decap_8 FILLER_20_977 ();
 sg13g2_decap_8 FILLER_20_984 ();
 sg13g2_decap_8 FILLER_20_991 ();
 sg13g2_decap_8 FILLER_20_998 ();
 sg13g2_decap_8 FILLER_20_1005 ();
 sg13g2_decap_8 FILLER_20_1012 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_21_424 ();
 sg13g2_decap_8 FILLER_21_431 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_decap_8 FILLER_21_445 ();
 sg13g2_decap_8 FILLER_21_452 ();
 sg13g2_decap_8 FILLER_21_459 ();
 sg13g2_decap_8 FILLER_21_466 ();
 sg13g2_decap_8 FILLER_21_473 ();
 sg13g2_decap_8 FILLER_21_480 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_8 FILLER_21_494 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_decap_8 FILLER_21_508 ();
 sg13g2_decap_8 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_522 ();
 sg13g2_decap_8 FILLER_21_529 ();
 sg13g2_decap_8 FILLER_21_536 ();
 sg13g2_decap_8 FILLER_21_543 ();
 sg13g2_decap_8 FILLER_21_550 ();
 sg13g2_decap_8 FILLER_21_557 ();
 sg13g2_decap_8 FILLER_21_564 ();
 sg13g2_decap_8 FILLER_21_571 ();
 sg13g2_decap_8 FILLER_21_578 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_592 ();
 sg13g2_decap_8 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_606 ();
 sg13g2_decap_8 FILLER_21_613 ();
 sg13g2_decap_8 FILLER_21_620 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_decap_8 FILLER_21_634 ();
 sg13g2_decap_8 FILLER_21_641 ();
 sg13g2_decap_8 FILLER_21_648 ();
 sg13g2_decap_8 FILLER_21_655 ();
 sg13g2_decap_8 FILLER_21_662 ();
 sg13g2_decap_8 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_676 ();
 sg13g2_decap_8 FILLER_21_683 ();
 sg13g2_decap_8 FILLER_21_690 ();
 sg13g2_decap_8 FILLER_21_697 ();
 sg13g2_decap_8 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_732 ();
 sg13g2_decap_8 FILLER_21_739 ();
 sg13g2_decap_8 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_753 ();
 sg13g2_decap_8 FILLER_21_760 ();
 sg13g2_decap_8 FILLER_21_767 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_decap_8 FILLER_21_781 ();
 sg13g2_decap_8 FILLER_21_788 ();
 sg13g2_decap_8 FILLER_21_795 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_decap_8 FILLER_21_809 ();
 sg13g2_decap_8 FILLER_21_816 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_decap_8 FILLER_21_837 ();
 sg13g2_decap_8 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_851 ();
 sg13g2_decap_8 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_21_865 ();
 sg13g2_decap_8 FILLER_21_872 ();
 sg13g2_decap_8 FILLER_21_879 ();
 sg13g2_decap_8 FILLER_21_886 ();
 sg13g2_decap_8 FILLER_21_893 ();
 sg13g2_decap_8 FILLER_21_900 ();
 sg13g2_decap_8 FILLER_21_907 ();
 sg13g2_decap_8 FILLER_21_914 ();
 sg13g2_decap_8 FILLER_21_921 ();
 sg13g2_decap_8 FILLER_21_928 ();
 sg13g2_decap_8 FILLER_21_935 ();
 sg13g2_decap_8 FILLER_21_942 ();
 sg13g2_decap_8 FILLER_21_949 ();
 sg13g2_decap_8 FILLER_21_956 ();
 sg13g2_decap_8 FILLER_21_963 ();
 sg13g2_decap_8 FILLER_21_970 ();
 sg13g2_decap_8 FILLER_21_977 ();
 sg13g2_decap_8 FILLER_21_984 ();
 sg13g2_decap_8 FILLER_21_991 ();
 sg13g2_decap_8 FILLER_21_998 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_fill_2 FILLER_21_1026 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_508 ();
 sg13g2_decap_8 FILLER_22_515 ();
 sg13g2_decap_8 FILLER_22_522 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_decap_8 FILLER_22_921 ();
 sg13g2_decap_8 FILLER_22_928 ();
 sg13g2_decap_8 FILLER_22_935 ();
 sg13g2_decap_8 FILLER_22_942 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_956 ();
 sg13g2_decap_8 FILLER_22_963 ();
 sg13g2_decap_8 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_decap_8 FILLER_22_991 ();
 sg13g2_decap_8 FILLER_22_998 ();
 sg13g2_decap_8 FILLER_22_1005 ();
 sg13g2_decap_8 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1019 ();
 sg13g2_fill_2 FILLER_22_1026 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_529 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_599 ();
 sg13g2_decap_8 FILLER_23_606 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_decap_8 FILLER_23_725 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_753 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_893 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_decap_8 FILLER_23_907 ();
 sg13g2_decap_8 FILLER_23_914 ();
 sg13g2_decap_8 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_935 ();
 sg13g2_decap_8 FILLER_23_942 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_963 ();
 sg13g2_decap_8 FILLER_23_970 ();
 sg13g2_decap_8 FILLER_23_977 ();
 sg13g2_decap_8 FILLER_23_984 ();
 sg13g2_decap_8 FILLER_23_991 ();
 sg13g2_decap_8 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_decap_8 FILLER_23_1012 ();
 sg13g2_decap_8 FILLER_23_1019 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_543 ();
 sg13g2_decap_8 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_620 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_879 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_decap_8 FILLER_24_907 ();
 sg13g2_decap_8 FILLER_24_914 ();
 sg13g2_decap_8 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_928 ();
 sg13g2_decap_8 FILLER_24_935 ();
 sg13g2_decap_8 FILLER_24_942 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_decap_8 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_445 ();
 sg13g2_decap_8 FILLER_25_452 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_8 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_494 ();
 sg13g2_decap_8 FILLER_25_501 ();
 sg13g2_decap_8 FILLER_25_508 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_decap_8 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_decap_8 FILLER_25_571 ();
 sg13g2_decap_8 FILLER_25_578 ();
 sg13g2_decap_8 FILLER_25_585 ();
 sg13g2_decap_8 FILLER_25_592 ();
 sg13g2_decap_8 FILLER_25_599 ();
 sg13g2_decap_8 FILLER_25_606 ();
 sg13g2_decap_8 FILLER_25_613 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_decap_8 FILLER_25_627 ();
 sg13g2_decap_8 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_641 ();
 sg13g2_decap_8 FILLER_25_648 ();
 sg13g2_decap_8 FILLER_25_655 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_25_865 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_decap_8 FILLER_25_893 ();
 sg13g2_decap_8 FILLER_25_900 ();
 sg13g2_decap_8 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_914 ();
 sg13g2_decap_8 FILLER_25_921 ();
 sg13g2_decap_8 FILLER_25_928 ();
 sg13g2_decap_8 FILLER_25_935 ();
 sg13g2_decap_8 FILLER_25_942 ();
 sg13g2_decap_8 FILLER_25_949 ();
 sg13g2_decap_8 FILLER_25_956 ();
 sg13g2_decap_8 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_970 ();
 sg13g2_decap_8 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_984 ();
 sg13g2_decap_8 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_998 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_8 FILLER_25_1012 ();
 sg13g2_decap_8 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_431 ();
 sg13g2_decap_8 FILLER_26_438 ();
 sg13g2_decap_8 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_decap_8 FILLER_26_466 ();
 sg13g2_decap_8 FILLER_26_473 ();
 sg13g2_decap_8 FILLER_26_480 ();
 sg13g2_decap_8 FILLER_26_487 ();
 sg13g2_decap_8 FILLER_26_494 ();
 sg13g2_decap_8 FILLER_26_501 ();
 sg13g2_decap_8 FILLER_26_508 ();
 sg13g2_decap_8 FILLER_26_515 ();
 sg13g2_decap_8 FILLER_26_522 ();
 sg13g2_decap_8 FILLER_26_529 ();
 sg13g2_decap_8 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_543 ();
 sg13g2_decap_8 FILLER_26_550 ();
 sg13g2_decap_8 FILLER_26_557 ();
 sg13g2_decap_8 FILLER_26_564 ();
 sg13g2_decap_8 FILLER_26_571 ();
 sg13g2_decap_8 FILLER_26_578 ();
 sg13g2_decap_8 FILLER_26_585 ();
 sg13g2_decap_8 FILLER_26_592 ();
 sg13g2_decap_8 FILLER_26_599 ();
 sg13g2_decap_8 FILLER_26_606 ();
 sg13g2_decap_8 FILLER_26_613 ();
 sg13g2_decap_8 FILLER_26_620 ();
 sg13g2_decap_8 FILLER_26_627 ();
 sg13g2_decap_8 FILLER_26_634 ();
 sg13g2_decap_8 FILLER_26_641 ();
 sg13g2_decap_8 FILLER_26_648 ();
 sg13g2_decap_8 FILLER_26_655 ();
 sg13g2_decap_8 FILLER_26_662 ();
 sg13g2_decap_8 FILLER_26_669 ();
 sg13g2_decap_8 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_683 ();
 sg13g2_decap_8 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_decap_8 FILLER_26_704 ();
 sg13g2_decap_8 FILLER_26_711 ();
 sg13g2_decap_8 FILLER_26_718 ();
 sg13g2_decap_8 FILLER_26_725 ();
 sg13g2_decap_8 FILLER_26_732 ();
 sg13g2_decap_8 FILLER_26_739 ();
 sg13g2_decap_8 FILLER_26_746 ();
 sg13g2_decap_8 FILLER_26_753 ();
 sg13g2_decap_8 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_781 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_8 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_26_865 ();
 sg13g2_decap_8 FILLER_26_872 ();
 sg13g2_decap_8 FILLER_26_879 ();
 sg13g2_decap_8 FILLER_26_886 ();
 sg13g2_decap_8 FILLER_26_893 ();
 sg13g2_decap_8 FILLER_26_900 ();
 sg13g2_decap_8 FILLER_26_907 ();
 sg13g2_decap_8 FILLER_26_914 ();
 sg13g2_decap_8 FILLER_26_921 ();
 sg13g2_decap_8 FILLER_26_928 ();
 sg13g2_decap_8 FILLER_26_935 ();
 sg13g2_decap_8 FILLER_26_942 ();
 sg13g2_decap_8 FILLER_26_949 ();
 sg13g2_decap_8 FILLER_26_956 ();
 sg13g2_decap_8 FILLER_26_963 ();
 sg13g2_decap_8 FILLER_26_970 ();
 sg13g2_decap_8 FILLER_26_977 ();
 sg13g2_decap_8 FILLER_26_984 ();
 sg13g2_decap_8 FILLER_26_991 ();
 sg13g2_decap_8 FILLER_26_998 ();
 sg13g2_decap_8 FILLER_26_1005 ();
 sg13g2_decap_8 FILLER_26_1012 ();
 sg13g2_decap_8 FILLER_26_1019 ();
 sg13g2_fill_2 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_decap_8 FILLER_28_431 ();
 sg13g2_decap_8 FILLER_28_438 ();
 sg13g2_decap_8 FILLER_28_445 ();
 sg13g2_decap_8 FILLER_28_452 ();
 sg13g2_decap_8 FILLER_28_459 ();
 sg13g2_decap_8 FILLER_28_466 ();
 sg13g2_decap_8 FILLER_28_473 ();
 sg13g2_decap_8 FILLER_28_480 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_8 FILLER_28_494 ();
 sg13g2_decap_8 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_508 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_522 ();
 sg13g2_decap_8 FILLER_28_529 ();
 sg13g2_decap_8 FILLER_28_536 ();
 sg13g2_decap_8 FILLER_28_543 ();
 sg13g2_decap_8 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_557 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_decap_8 FILLER_28_571 ();
 sg13g2_decap_8 FILLER_28_578 ();
 sg13g2_decap_8 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_8 FILLER_28_606 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_8 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_956 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_fill_2 FILLER_28_1026 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_decap_8 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_882 ();
 sg13g2_decap_8 FILLER_29_889 ();
 sg13g2_decap_8 FILLER_29_896 ();
 sg13g2_decap_8 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_910 ();
 sg13g2_decap_8 FILLER_29_917 ();
 sg13g2_decap_8 FILLER_29_924 ();
 sg13g2_decap_8 FILLER_29_931 ();
 sg13g2_decap_8 FILLER_29_938 ();
 sg13g2_decap_8 FILLER_29_945 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_decap_8 FILLER_29_959 ();
 sg13g2_decap_8 FILLER_29_966 ();
 sg13g2_decap_8 FILLER_29_973 ();
 sg13g2_decap_8 FILLER_29_980 ();
 sg13g2_decap_8 FILLER_29_987 ();
 sg13g2_decap_8 FILLER_29_994 ();
 sg13g2_decap_8 FILLER_29_1001 ();
 sg13g2_decap_8 FILLER_29_1008 ();
 sg13g2_decap_8 FILLER_29_1015 ();
 sg13g2_decap_8 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_decap_8 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_938 ();
 sg13g2_decap_8 FILLER_32_945 ();
 sg13g2_decap_8 FILLER_32_952 ();
 sg13g2_decap_8 FILLER_32_959 ();
 sg13g2_decap_8 FILLER_32_966 ();
 sg13g2_decap_8 FILLER_32_973 ();
 sg13g2_decap_8 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_8 FILLER_34_896 ();
 sg13g2_decap_8 FILLER_34_903 ();
 sg13g2_decap_8 FILLER_34_910 ();
 sg13g2_decap_8 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_decap_8 FILLER_35_875 ();
 sg13g2_decap_8 FILLER_35_882 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_decap_8 FILLER_35_896 ();
 sg13g2_decap_8 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_910 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_945 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_8 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_973 ();
 sg13g2_decap_8 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_8 FILLER_35_994 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_36_868 ();
 sg13g2_decap_8 FILLER_36_875 ();
 sg13g2_decap_8 FILLER_36_882 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_decap_8 FILLER_36_896 ();
 sg13g2_decap_8 FILLER_36_903 ();
 sg13g2_decap_8 FILLER_36_910 ();
 sg13g2_decap_8 FILLER_36_917 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_decap_8 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_39_931 ();
 sg13g2_decap_8 FILLER_39_938 ();
 sg13g2_decap_8 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_966 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_decap_8 FILLER_39_980 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_40_868 ();
 sg13g2_decap_8 FILLER_40_875 ();
 sg13g2_decap_8 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_889 ();
 sg13g2_decap_8 FILLER_40_896 ();
 sg13g2_decap_8 FILLER_40_903 ();
 sg13g2_decap_8 FILLER_40_910 ();
 sg13g2_decap_8 FILLER_40_917 ();
 sg13g2_decap_8 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_decap_8 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_8 FILLER_41_917 ();
 sg13g2_decap_8 FILLER_41_924 ();
 sg13g2_decap_8 FILLER_41_931 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_8 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_994 ();
 sg13g2_decap_8 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_decap_8 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_882 ();
 sg13g2_decap_8 FILLER_42_889 ();
 sg13g2_decap_8 FILLER_42_896 ();
 sg13g2_decap_8 FILLER_42_903 ();
 sg13g2_decap_8 FILLER_42_910 ();
 sg13g2_decap_8 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_924 ();
 sg13g2_decap_8 FILLER_42_931 ();
 sg13g2_decap_8 FILLER_42_938 ();
 sg13g2_decap_8 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_966 ();
 sg13g2_decap_8 FILLER_42_973 ();
 sg13g2_decap_8 FILLER_42_980 ();
 sg13g2_decap_8 FILLER_42_987 ();
 sg13g2_decap_8 FILLER_42_994 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_532 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_875 ();
 sg13g2_decap_8 FILLER_44_882 ();
 sg13g2_decap_8 FILLER_44_889 ();
 sg13g2_decap_8 FILLER_44_896 ();
 sg13g2_decap_8 FILLER_44_903 ();
 sg13g2_decap_8 FILLER_44_910 ();
 sg13g2_decap_8 FILLER_44_917 ();
 sg13g2_decap_8 FILLER_44_924 ();
 sg13g2_decap_8 FILLER_44_931 ();
 sg13g2_decap_8 FILLER_44_938 ();
 sg13g2_decap_8 FILLER_44_945 ();
 sg13g2_decap_8 FILLER_44_952 ();
 sg13g2_decap_8 FILLER_44_959 ();
 sg13g2_decap_8 FILLER_44_966 ();
 sg13g2_decap_8 FILLER_44_973 ();
 sg13g2_decap_8 FILLER_44_980 ();
 sg13g2_decap_8 FILLER_44_987 ();
 sg13g2_decap_8 FILLER_44_994 ();
 sg13g2_decap_8 FILLER_44_1001 ();
 sg13g2_decap_8 FILLER_44_1008 ();
 sg13g2_decap_8 FILLER_44_1015 ();
 sg13g2_decap_8 FILLER_44_1022 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_decap_8 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_decap_8 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_decap_8 FILLER_45_952 ();
 sg13g2_decap_8 FILLER_45_959 ();
 sg13g2_decap_8 FILLER_45_966 ();
 sg13g2_decap_8 FILLER_45_973 ();
 sg13g2_decap_8 FILLER_45_980 ();
 sg13g2_decap_8 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net;
 assign uio_out[3] = net1;
 assign uio_out[4] = net2;
 assign uio_out[5] = net3;
 assign uio_out[6] = net4;
 assign uio_out[7] = net5;
 assign uo_out[0] = net6;
 assign uo_out[1] = net7;
 assign uo_out[2] = net8;
 assign uo_out[3] = net9;
 assign uo_out[4] = net10;
 assign uo_out[5] = net11;
 assign uo_out[6] = net12;
 assign uo_out[7] = net13;
endmodule
